��      �Player�h ��)��}�(�char��@��armorPen�K �range�K�level�K�
hitEffects�]��leftRing�N�recalcTimer�K �expNext�K��skills�}�(�3��	Abilities��Fireball����2�h�Shocking_Grasp����7�h�Ready_for_Battle����4�h�Lightning_Bolt����6�h�Rending_Blow����5�h�Block����1�h�Charge���u�power�K�dodge�K �visible���	rightRing�N�canMove���	recalcMax�K �
countering���
prevTarget�N�skillPoints�K�leftHand��Items.Weapons��Tome���)��}�(�
consumable��h&K �weight�K�type��0H��addPower��hK�name�h1�
usesArrows��hKh�?��color�]�(K�K�K�e�	throwable���
equippable��hK �magPower�Kub�health�K1�blocking���
leftScroll�N�arrows�K�	rightHand�h0�
Greatsword���)��}�(h5�h&Kh6Kh7�2H�h9�hKh:hGh;�hKhh<h=h>h?�h@�hKhAKub�invertColor���
initiative�K�gold�MS�items�]�(�Items.Armors��Leather_Helm���)��}�(h6KhKh7�helmet��pObject�Nh=h>h?�h@�h5��armorVal�K
hh<h:�Leather Helm�ubhQ�Leather_Shirt���)��}�(h6KhKh7�armor�hWNh=h>h?�h@�h5�hXKhh<h:�Leather Shirt�ubh[)��}�(h6KhKh7h^hWNh=h>h?�h@�h5�hXKhh<h:h_ubh0�Spear���)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hbh;�hKhh<h=h>h?�h@�hKhAKubhQ�	Iron_Helm���)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:�	Iron Helm�ubh0�	Longsword���)��}�(hWNh5�h&Kh6Kh7�1H�h9�hKh:hkh;�hKhh<h=h>h?�h@�hKhAKubh[)��}�(h6KhKh7h^hWNh=h>h?�h@�h5�hXKhh<h:h_ubh0�Wooden_Shield���)��}�(hWNh5�h&K h6KhXKh7hoh9�hKh:�Wooden Shield�h;�hKhh<h=h>h?�h@�hAK ubhQ�	Cloth_Hat���)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:�	Cloth Hat�ubhx)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:h{ubhQ�Chain_Shirt���)��}�(h6K#hKh7h^h=h>h?�h@�h5�hXK#hh<h:�Chain Shirt�ub�Items.Consumables��Scroll_of_Fireball���)��}�(hWNhKh7�scroll�h=h>h@�h5�h�s��spell�hh:�Scroll of Fireball�ubhg)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:hjubhx)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:h{ubhx)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:h{ubh0�Bow���)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubh�)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhl)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:hkh;�hKhh<h=h>h?�h@�hKhAKubhl)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:hkh;�hKhh<h=h>h?�h@�hKhAKubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubh[)��}�(h6KhKh7h^hWNh=h>h?�h@�h5�hXKhh<h:h_ubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhH)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hGh;�hKhh<h=h>h?�h@�hKhAKubhg)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:hjubh[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhH)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hGh;�hKhh<h=h>h?�h@�hKhAKubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubh�)��}�(hWNhKh7h�h=h>h@�h5�hh�h�hh:h�ubhc)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hbh;�hKhh<h=h>h?�h@�hKhAKubhx)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:h{ubh�)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubh[)��}�(h6KhKh7h^hWNh=h>h?�h@�h5�hXKhh<h:h_ubhs)��}�(hWNh5�h&K h6KhXKh7hoh9�hKh:hvh;�hKhh<h=h>h?�h@�hAK ubh[)��}�(h6KhKh7h^hWNh=h>h?�h@�h5�hXKhh<h:h_ubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhg)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:hjubhx)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:h{ubhg)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:hjubh�)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubh0�Mace���)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubh�)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhc)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hbh;�hKhh<h=h>h?�h@�hKhAKubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubh0�Dagger���)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhH)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hGh;�hKhh<h=h>h?�h@�hKhAKubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhx)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:h{ubhQ�Cloth_Shirt���)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:�Cloth Shirt�ubhc)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hbh;�hKhh<h=h>h?�h@�hKhAKubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhx)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:h{ubh�)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhl)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:hkh;�hKhh<h=h>h?�h@�hKhAKubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhl)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:hkh;�hKhh<h=h>h?�h@�hKhAKubh)��}�(h6K#hKh7h^h=h>h?�h@�h5�hXK#hh<h:h�ubh��	Time_Bomb���)��}�(h5��radius�Kh7h5hK h:�Bomb��dur�KhKh�o�h=h>�damage�Kh@��desc��Explodes up after 3 turns�ubhQ�
Chain_Helm���)��}�(h6K
hKh7hVh=h>h?�h@�h5�hXKhh<h:�
Chain Helm�ubhx)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:h{ubh�)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhx)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:h{ubhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYubhx)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:h{ubhx)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:h{ubh�)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubh0�Iron_Shield���)��}�(hWNh5�h&K h6KhXKh7hoh9�hKh:�Iron Shield�h;�hKhh<h=h>h?�h@�hAK ubhx)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:h{ubh�)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubh[)��}�(h6KhKh7h^hWNh=h>h?�h@�h5�hXKhh<h:h_ubh�)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhg)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:hjubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhl)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:hkh;�hKhh<h=h>h?�h@�hKhAKubh�)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhH)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hGh;�hKhh<h=h>h?�h@�hKhAKubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubh�)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhc)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hbh;�hKhh<h=h>h?�h@�hKhAKubhc)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hbh;�hKhh<h=h>h?�h@�hKhAKubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhx)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:h{ubhc)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hbh;�hKhh<h=h>h?�h@�hKhAKubh�)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubh�)��}�(hWNh5�h�Kh7h5hK h:h�h�KhKhh�h=h>h�Kh@�h�h�ubhx)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:h{ubh�)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubh�)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h�ubh�)��}�(hKh7h�h=h>h@�h5�hh�h�hh:h�ubhs)��}�(h5�h&K h6KhXKh7hoh9�hKh:hvh;�hKhh<h=h>h?�h@�hAK ubh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhg)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:hjubh�)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h�ubh�)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubh�)��}�(hWNhKh7h�h=h>h@�h5�hh�h�hh:h�ubh[)��}�(h6KhKh7h^hWNh=h>h?�h@�h5�hXKhh<h:h_ubhg)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:hjubh[)��}�(h6KhKh7h^hWNh=h>h?�h@�h5�hXKhh<h:h_ubhl)��}�(h5�h&Kh6Kh7hoh9�hKh:hkh;�hKhh<h=h>h?�h@�hKhAKubh�)��}�(h5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhc)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hbh;�hKhh<h=h>h?�h@�hKhAKubh��	GreenHerb���)��}�(hWNh7h5h=h>h@�h5�h�+��healNum�Kh:�
Green Herb�ubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhS)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXK
hh<h:hYubhH)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hGh;�hKhh<h=h>h?�h@�hKhAKubh[)��}�(h6KhKh7h^hWNh=h>h?�h@�h5�hXKhh<h:h_ubhH)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hGh;�hKhh<h=h>h?�h@�hKhAKubh�)��}�(hWNh5�h�Kh7h5hK h:h�h�KhKhh�h=h>h�Kh@�h�h�ubh�)��}�(hWNh5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhg)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:hjubh�)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKube�exp�K��
baseHealth�M�
healthTemp�K �effects�]�hXK �	healthMax�M,�playerControlled���skillLevels�}�(hKhKhK hKhK h K h#K uh:�George�hW�Object�j�  ��)��}�(�col�KE�pLevel��LevelTypes.LevelTypes��Tower���)��}�(�	thePlayer�h�levelManager��LevelManager�j�  ��)��}�(�cursor�K �	levelList�]�j�  a�
messageSys��
MessageSys��Messages���)��}�(�retrieveLimit�K�messageLimit�M��messages�]�(�Goblin Grunt dropped Longsword��!Goblin Grunt dropped Leather Helm��Goblin Grunt dropped Buckler��!Goblin Grunt was killed by George��Goblin Grunt is afraid!��"George attacked Goblin Grunt for 4��Goblin Grunt missed George��George acquired 5 coins��"Goblin Grunt attacked George for 3��George picked up Bow�� Goblin Grunt picked up Cloth Hat�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 4��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George picked up Iron Helm��#Goblin Archer attacked George for 1��#Goblin Berserker dropped Gold Coins��&Goblin Berserker dropped Leather Shirt��"Goblin Berserker dropped Iron Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 4��#Goblin Archer attacked George for 1��&Goblin Berserker attacked George for 5��George acquired 12 coins��#Goblin Archer attacked George for 1��&Goblin Berserker attacked George for 5��George picked up Mace��#Goblin Archer attacked George for 1��$Goblin Berserker picked up Iron Helm��#Goblin Stonewall dropped Gold Coins��Goblin Stonewall dropped Mace��"Goblin Stonewall dropped Iron Helm��%Goblin Stonewall was killed by George��Goblin Stonewall is afraid!��&George attacked Goblin Stonewall for 2��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��&George attacked Goblin Berserker for 2��&George attacked Goblin Stonewall for 2��George used Fireball��&Goblin Stonewall attacked George for 3��&George attacked Goblin Berserker for 2��&George attacked Goblin Stonewall for 2��George used Lightning Bolt��George waited...��George waited...��George waited...��George picked up Bomb��George picked up Greatsword��George picked up Leather Shirt��George picked up Greatsword��George picked up Leather Helm��#Goblin Berserker dropped Greatsword��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 4��&Goblin Berserker attacked George for 5��&George attacked Goblin Berserker for 4��&Goblin Berserker attacked George for 5��George picked up Leather Helm��#Goblin Berserker dropped Greatsword��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 4��&Goblin Berserker attacked George for 5��George picked up Leather Helm��Goblin Berserker dropped Bomb��&Goblin Berserker dropped Leather Shirt��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 4��&Goblin Berserker attacked George for 5��George picked up Green Herb��&Goblin Berserker attacked George for 5��George picked up Spear��'Goblin Berserker picked up Leather Helm�� Goblin Lancer dropped Green Herb��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 4��Goblin Lancer missed George��#Goblin Lancer attacked George for 2��&George attacked Goblin Berserker for 2��&George attacked Goblin Berserker for 2��George used Fireball��#Goblin Lancer attacked George for 2��&George attacked Goblin Berserker for 2��#George attacked Goblin Lancer for 2��George used Lightning Bolt��George waited...��George waited...��George waited...��George acquired 8 coins��George picked up Bow��George acquired 8 coins��George picked up Longsword��George acquired 9 coins��George picked up Leather Shirt��George picked up Iron Helm��#Goblin Berserker dropped Gold Coins��&Goblin Berserker dropped Leather Shirt��"Goblin Berserker dropped Iron Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 4��&Goblin Berserker attacked George for 5��George acquired 5 coins��&Goblin Berserker attacked George for 5��George picked up Leather Shirt��$Goblin Berserker picked up Iron Helm��Goblin Grunt dropped Gold Coins��"Goblin Grunt dropped Leather Shirt��Goblin Grunt dropped Iron Helm��!Goblin Grunt was killed by George��Goblin Grunt is afraid!��"George attacked Goblin Grunt for 4��Goblin Grunt missed George��#George picked up Scroll of Fireball��"Goblin Grunt attacked George for 3��George picked up Mace�� Goblin Grunt picked up Iron Helm��+Goblin Stonewall dropped Scroll of Fireball��Goblin Stonewall dropped Mace��"Goblin Stonewall dropped Iron Helm��%Goblin Stonewall was killed by George��Goblin Stonewall is afraid!��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&George attacked Goblin Stonewall for 2��"George attacked Goblin Grunt for 2��George used Fireball��&George attacked Goblin Berserker for 2��George missed Goblin Grunt��&George attacked Goblin Stonewall for 2��George used Lightning Bolt��George acquired 8 coins��George picked up Cloth Shirt��George picked up Iron Helm��George picked up Dagger��George acquired 12 coins��George picked up Wooden Shield��#George picked up Scroll of Fireball��George picked up Cloth Shirt��George picked up Bow��George picked up Cloth Hat��George acquired 10 coins��George picked up Bomb��George acquired 13 coins��George acquired 12 coins��George picked up Bow��George picked up Spear��George picked up Cloth Hat��George picked up Leather Helm��George picked up Spear��George picked up Spear�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 6��George used Shocking Grasp��George used Shocking Grasp�� Goblin Lancer dropped Gold Coins��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 4��#Goblin Lancer attacked George for 2��George picked up Leather Helm��#Goblin Lancer attacked George for 2��#George attacked Goblin Lancer for 2��George used Lightning Bolt��#Goblin Lancer attacked George for 2��Goblin Lancer dropped Bomb��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 4��#Goblin Lancer attacked George for 2��#Goblin Lancer attacked George for 2��George picked up Leather Helm�� Goblin Lancer dropped Gold Coins��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 4��#Goblin Lancer attacked George for 2��#Goblin Archer attacked George for 1��#Goblin Lancer attacked George for 2��#Goblin Archer attacked George for 1��George waited...��#Goblin Archer attacked George for 1��George waited...��#Goblin Archer attacked George for 1��George waited...��#Goblin Archer attacked George for 1�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 4��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George waited...��George acquired 5 coins��George picked up Dagger��George picked up Leather Helm��Goblin Thief dropped Gold Coins��Goblin Thief dropped Dagger��!Goblin Thief dropped Leather Helm��!Goblin Thief was killed by George��"George attacked Goblin Thief for 2��George used Lightning Bolt��George used a Green Herb��George used a Green Herb��George used a Green Herb��George acquired 11 coins��George acquired 4 coins��George picked up Greatsword��George picked up Mace��George picked up Longsword��George picked up Leather Helm��Goblin Grunt dropped Gold Coins��Goblin Grunt dropped Longsword��!Goblin Grunt dropped Leather Helm��!Goblin Grunt was killed by George��Goblin Grunt is afraid!��"George attacked Goblin Grunt for 4��"Goblin Grunt attacked George for 3��George picked up Iron Helm��#Goblin Stonewall dropped Gold Coins��Goblin Stonewall dropped Mace��"Goblin Stonewall dropped Iron Helm��%Goblin Stonewall was killed by George��Goblin Stonewall is afraid!��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��Goblin Stonewall missed George��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&Goblin Stonewall attacked George for 3��George picked up Leather Helm��&George attacked Goblin Stonewall for 2��#Goblin Berserker dropped Greatsword��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 2��George used Fireball��&Goblin Berserker attacked George for 5��&George attacked Goblin Stonewall for 2��&George attacked Goblin Berserker for 2��George used Lightning Bolt��George waited...��"George attacked Goblin Grunt for 2��George used Lightning Bolt��"George attacked Goblin Thief for 2��&George attacked Goblin Berserker for 2��George used Fireball��George acquired 6 Arrows��George picked up Dagger��George picked up Leather Shirt��George picked up Bow��George picked up Cloth Hat��George picked up Iron Shield��Goblin Thief dropped Dagger��"Goblin Thief dropped Leather Shirt�� Goblin Thief dropped Iron Shield��!Goblin Thief was killed by George��"George attacked Goblin Thief for 2��George used Lightning Bolt��&Goblin Archer dropped Bundle of Arrows��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��#George attacked Goblin Archer for 2��"George attacked Goblin Thief for 2��George used Fireball��George acquired 14 coins��George picked up Bow��George picked up Cloth Hat�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��#George attacked Goblin Archer for 4��#Goblin Archer attacked George for 1��George acquired 10 coins��George picked up Cloth Hat��George picked up Leather Helm��George picked up Cloth Hat��George picked up Bow��George picked up Cloth Hat��"Goblin Thief picked up Iron Shield��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 4��George acquired 16 coins��George picked up Chain Helm��George picked up Bomb��George picked up Chain Shirt��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George picked up Longsword��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George picked up Leather Helm��#Goblin Archer attacked George for 1��Goblin Grunt dropped Longsword��!Goblin Grunt dropped Leather Helm��!Goblin Grunt was killed by George��Goblin Grunt is afraid!��"George attacked Goblin Grunt for 4��"George attacked Goblin Grunt for 2��George used Lightning Bolt��George waited...��George picked up Longsword��George acquired 12 coins��George picked up Bow��George picked up Cloth Hat�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 6��George used Shocking Grasp��George used Shocking Grasp��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George picked up Leather Helm��#Goblin Archer attacked George for 1��Goblin Archer is afraid!��#George attacked Goblin Archer for 2��Goblin Grunt dropped Longsword��!Goblin Grunt dropped Leather Helm��!Goblin Grunt was killed by George��Goblin Grunt is afraid!��"George attacked Goblin Grunt for 2��George used Fireball��Goblin Archer is afraid!��#George attacked Goblin Archer for 2��"George attacked Goblin Grunt for 2��George used Lightning Bolt��#Goblin Archer attacked George for 1��George waited...��#Goblin Archer attacked George for 1��George acquired 8 coins��George picked up Spear��George acquired 10 coins��George acquired 7 Arrows��George picked up Cloth Shirt��George picked up Cloth Hat��George picked up Leather Helm�� Goblin Lancer dropped Gold Coins��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 4��#Goblin Lancer attacked George for 2��#Goblin Lancer attacked George for 2��George waited...��#Goblin Lancer attacked George for 2��George picked up Greatsword��George picked up Leather Helm��#Goblin Berserker dropped Greatsword��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 6��George used Shocking Grasp��George used Shocking Grasp��George missed Goblin Lancer��George used Lightning Bolt��George acquired 5 coins��George picked up Dagger��George picked up Leather Helm��Goblin Thief dropped Gold Coins��Goblin Thief dropped Dagger��!Goblin Thief dropped Leather Helm��!Goblin Thief was killed by George��"George attacked Goblin Thief for 4��"Goblin Thief attacked George for 3��George waited...��George waited...��George waited...��George acquired 12 coins��George acquired 7 Arrows��George acquired 12 coins��George picked up Spear��George picked up Mace��George picked up Mace��George picked up Bow��George picked up Iron Helm��George leveled up!��)Goblin Stonewall dropped Bundle of Arrows��Goblin Stonewall dropped Mace��"Goblin Stonewall dropped Iron Helm��%Goblin Stonewall was killed by George��Goblin Stonewall is afraid!��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��Goblin Stonewall missed George��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��George picked up Cloth Hat��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 3��#Goblin Archer attacked George for 1��George picked up Iron Helm��#Goblin Stonewall dropped Gold Coins��Goblin Stonewall dropped Mace��"Goblin Stonewall dropped Iron Helm��%Goblin Stonewall was killed by George��Goblin Stonewall is afraid!��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��George picked up Leather Helm�� Goblin Lancer dropped Gold Coins��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 3��#Goblin Lancer attacked George for 2��#George attacked Goblin Lancer for 3��#Goblin Lancer attacked George for 2��Goblin Lancer missed George��George acquired 7 coins��George picked up Leather Shirt��George picked up Wooden Shield��George acquired 5 coins��George picked up Leather Shirt��George picked up Bow��George picked up Cloth Hat�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 3��#Goblin Archer attacked George for 1��George picked up Spear��#Goblin Archer attacked George for 1��#Goblin Knight dropped Wooden Shield��#Goblin Knight dropped Leather Shirt��Goblin Knight dropped Spear��"Goblin Knight was killed by George��Goblin Knight is afraid!��#George attacked Goblin Knight for 3��#Goblin Knight attacked George for 4��#Goblin Archer attacked George for 1��#George attacked Goblin Knight for 3��#Goblin Knight attacked George for 4��#Goblin Archer attacked George for 1��George missed Goblin Knight��#Goblin Knight attacked George for 4��#Goblin Archer attacked George for 1��George missed Goblin Knight��Goblin Knight missed George��#Goblin Archer attacked George for 1��George missed Goblin Knight��#Goblin Knight attacked George for 4��#Goblin Archer attacked George for 1��#George picked up Scroll of Fireball��#Goblin Knight attacked George for 4��#Goblin Archer attacked George for 1��George picked up Leather Helm��#Goblin Knight attacked George for 4�� Goblin Archer dropped Gold Coins��#Goblin Archer dropped Leather Shirt��"Goblin Archer dropped Leather Helm��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 3��Goblin Knight picked up Spear��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George waited...��$Goblin Archer picked up Leather Helm��#Goblin Archer attacked George for 1��George picked up Greatsword��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George picked up Leather Helm��Goblin Archer missed George��#Goblin Archer attacked George for 1��#Goblin Berserker dropped Greatsword��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 3��#Goblin Archer attacked George for 1��&Goblin Berserker attacked George for 5��&George attacked Goblin Berserker for 3��#Goblin Archer attacked George for 1��&Goblin Berserker attacked George for 5��George missed Goblin Berserker��(Goblin Lancer dropped Scroll of Fireball��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 2��George used Lightning Bolt��&George attacked Goblin Berserker for 2��#George attacked Goblin Lancer for 2��George used Fireball��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George waited...��#Goblin Archer attacked George for 1��George acquired 11 coins��Goblin Archer missed George��George acquired 8 coins��George picked up Green Herb��George picked up Leather Shirt��George picked up Iron Helm��George acquired 11 coins��George picked up Greatsword��George waited...��George waited...��George acquired 8 coins��George picked up Leather Helm��#Goblin Berserker dropped Gold Coins��#Goblin Berserker dropped Greatsword��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 6��George used Shocking Grasp��George used Shocking Grasp��George picked up Leather Shirt��George picked up Leather Helm��#Goblin Berserker dropped Gold Coins��&Goblin Berserker dropped Leather Shirt��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 3��&Goblin Berserker attacked George for 5��George picked up Longsword��'Goblin Berserker picked up Leather Helm��George waited...��&George attacked Goblin Berserker for 2��Goblin Grunt dropped Longsword��!Goblin Grunt dropped Leather Helm��!Goblin Grunt was killed by George��Goblin Grunt is afraid!��"George attacked Goblin Grunt for 2��George used Fireball��"Goblin Grunt attacked George for 3��&George attacked Goblin Berserker for 2��"George attacked Goblin Grunt for 2��George used Lightning Bolt��George waited...��George waited...��George acquired 5 Arrows��George picked up Longsword��George acquired 6 coins��George acquired 4 coins��George picked up Bow��George picked up Bow��George picked up Cloth Hat�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 3��#Goblin Archer attacked George for 1��George picked up Cloth Hat��#Goblin Archer attacked George for 1�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 3��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George missed Goblin Archer��Goblin Archer missed George��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George picked up Iron Helm��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��&Goblin Knight dropped Bundle of Arrows��Goblin Knight dropped Longsword��Goblin Knight dropped Iron Helm��"Goblin Knight was killed by George��Goblin Knight is afraid!��#George attacked Goblin Knight for 3��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Knight attacked George for 4��#George attacked Goblin Knight for 3��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#George picked up Scroll of Fireball��George acquired 15 coins��George picked up Chain Shirt��George picked up Cloth Hat��George acquired 12 coins��George picked up Cloth Hat��George picked up Wooden Shield��George acquired 6 coins��George picked up Leather Shirt��George picked up Longsword��George picked up Iron Helm�� Goblin Knight dropped Gold Coins��Goblin Knight dropped Longsword��Goblin Knight dropped Iron Helm��"Goblin Knight was killed by George��Goblin Knight is afraid!��#George attacked Goblin Knight for 3��#Goblin Knight attacked George for 4��George picked up Spear��#Goblin Knight dropped Wooden Shield��#Goblin Knight dropped Leather Shirt��Goblin Knight dropped Spear��"Goblin Knight was killed by George��Goblin Knight is afraid!��#George attacked Goblin Knight for 3��#Goblin Knight attacked George for 4��#George attacked Goblin Knight for 3��#Goblin Knight attacked George for 4��George acquired 6 Arrows��#Goblin Knight attacked George for 4��George picked up Leather Shirt��Goblin Knight picked up Spear��)Goblin Berserker dropped Bundle of Arrows��&Goblin Berserker dropped Leather Shirt��Goblin Berserker dropped Spear��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 3��&Goblin Berserker attacked George for 5��George acquired 12 coins��&Goblin Berserker attacked George for 5��George picked up Leather Shirt��Goblin Berserker missed George��George picked up Leather Helm��&Goblin Berserker attacked George for 5��&George attacked Goblin Berserker for 2��#George attacked Goblin Knight for 2��#George attacked Goblin Knight for 2��George used Fireball��&Goblin Berserker attacked George for 5��George acquired 13 coins�� Goblin Berserker picked up Spear��George waited...��#Goblin Berserker dropped Gold Coins��&Goblin Berserker dropped Leather Shirt��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 6��George used Shocking Grasp��George used Shocking Grasp��'Goblin Berserker picked up Leather Helm��&George attacked Goblin Berserker for 2��#George attacked Goblin Knight for 2��&George attacked Goblin Berserker for 2�� Goblin Lancer dropped Gold Coins��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 2��George used Lightning Bolt��#Goblin Lancer attacked George for 2��#Goblin Lancer attacked George for 2��George waited...��George waited...��#George attacked Goblin Lancer for 2��&George attacked Goblin Berserker for 2��George used Fireball��Player Ready: George��
Game Start�eub�	gameState��__main__��Game���)��}�(�loadRequest��j�  h�width�K#�turn�M{	j�  j�  �xConst�K�yConst�KF�MessageHandler�j�  �height�K�console��tdl��Console���)��K_K/]�(K K K K ��K K K ����KGK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KLK�K�K���K K K ����KEK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KRK�K�K���K K K ����KPK�K�K���K K K ����KAK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KWK�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KxK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KaK�K�K���K K K ����KoK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KFK�K�K���K K K ����K K K K ��K K K ����KvK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KnK�K�K���K K K ����KwK�K�K���K K K ����KmK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KoK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KoK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KoK�K�K���K K K ����KbK�K�K���K K K ����KoK�K�K���K K K ����KbK�K�K���K K K ����KoK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KwK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KgK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KgK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KgK�K�K���K K K ����KiK�K�K���K K K ����KgK�K�K���K K K ����KiK�K�K���K K K ����KgK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K1K�K�K���K K K ����K K K K ��K K K ����KhK�K�K���K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K:K�K�K���K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KPK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K1K�K�K���K K K ����K5K�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KpK�K�K���K K K ����KAK�K�K���K K K ����KAK�K�K���K K K ����KaK�K�K���K K K ����KAK�K�K���K K K ����KAK�K�K���K K K ����KAK�K�K���K K K ����KAK�K�K���K K K ����KAK�K�K���K K K ����KGK�K�K���K K K ����KpK�K�K���K K K ����KGK�K�K���K K K ����KaK�K�K���K K K ����KGK�K�K���K K K ����KaK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K4K�K�K���K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K9K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KiK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KtK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KiK�K�K���K K K ����KrK�K�K���K K K ����KcK�K�K���K K K ����KrK�K�K���K K K ����KtK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KAK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K9K�K�K���K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KtK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KuK�K�K���K K K ����KcK�K�K���K K K ����KuK�K�K���K K K ����KqK�K�K���K K K ����KuK�K�K���K K K ����KtK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K9K�K�K���K K K ����K K K K ��K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KkK�K�K���K K K ����KhK�K�K���K K K ����KhK�K�K���K K K ����KaK�K�K���K K K ����KhK�K�K���K K K ����KhK�K�K���K K K ����KhK�K�K���K K K ����KhK�K�K���K K K ����KhK�K�K���K K K ����KnK�K�K���K K K ����KkK�K�K���K K K ����KnK�K�K���K K K ����KuK�K�K���K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KcK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KtK�K�K���K K K ����KeK�K�K���K K K ����KtK�K�K���K K K ����KiK�K�K���K K K ����KtK�K�K���K K K ����KcK�K�K���K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KSK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KdK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KkK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K�K�K���K K K ����KdK�K�K���K K K ����K K�K�K���K K K ����KrK�K�K���K K K ����K K�K�K���K K K ����KkK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KpK�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����KmK�K�K���K K K ����KeK�K�K���K K K ����KiK�K�K���K K K ����KwK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KcK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KuK�K�K���K K K ����KaK�K�K���K K K ����KaK�K�K���K K K ����KdK�K�K���K K K ����KiK�K�K���K K K ����KwK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KiK�K�K���K K K ����KuK�K�K���K K K ����KtK�K�K���K K K ����KdK�K�K���K K K ����KiK�K�K���K K K ����KdK�K�K���K K K ����KsK�K�K���K K K ����KaK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KkK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KpK�K�K���K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����KaK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KcK�K�K���K K K ����KpK�K�K���K K K ����KtK�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����KGK�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KkK�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����K5K�K�K���K K K ����KsK�K�K���K K K ����KGK�K�K���K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KIK�K�K���K K K ����KaK�K�K���K K K ����KaK�K�K���K K K ����KoK�K�K���K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KeK�K�K���K K K ����KBK�K�K���K K K ����KcK�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����KfK�K�K���K K K ����KkK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KrK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KbK�K�K���K K K ����KfK�K�K���K K K ����KkK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KdK�K�K���K K K ����KoK�K�K���K K K ����KkK�K�K���K K K ����KcK�K�K���K K K ����KdK�K�K���K K K ����KbK�K�K���K K K ����KrK�K�K���K K K ����KiK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KTK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KoK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KlK�K�K���K K K ����KrK�K�K���K K K ����KiK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����KwK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����KlK�K�K���K K K ����KaK�K�K���K K K ����KlK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KiK�K�K���K K K ����KaK�K�K���K K K ����KlK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KuK�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����KiK�K�K���K K K ����KGK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KwK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KnK�K�K���K K K ����KiK�K�K���K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����KnK�K�K���K K K ����KdK�K�K���K K K ����KeK�K�K���K K K ����KBK�K�K���K K K ����KLK�K�K���K K K ����KLK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KHK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KdK�K�K���K K K ����KeK�K�K���K K K ����KCK�K�K���K K K ����KBK�K�K���K K K ����KGK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����KsK�K�K���K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����K!K�K�K���K K K ����KdK�K�K���K K K ����KuK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KAK�K�K���K K K ����K!K�K�K���K K K ����KdK�K�K���K K K ����KlK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KCK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KcK�K�K���K K K ����KaK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KlK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KoK�K�K���K K K ����KwK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KbK�K�K���K K K ����KkK�K�K���K K K ����KtK�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KmK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KcK�K�K���K K K ����K K K K ��K K K ����KbK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KuK�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����KlK�K�K���K K K ����KhK�K�K���K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KwK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KgK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KCK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KrK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KfK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KfK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����KdK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����KfK�K�K���K K K ����KfK�K�K���K K K ����KfK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KsK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K �      K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K4K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K1K�K�K���K K K ����K4K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����e(K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K$K�K�K��K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K@KKYK���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K?K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K=KQKOK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K4K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KSK�K�K���K K K ����KLK�K�K���K K K ����KRK�K�K���K K K ����KDK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KFK�K�K���K K K ����KLK�K�K���K K K ����KRK�K�K���K K K ����KDK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KLK�K�K���K K K ����KLK�K�K���K K K ����KRK�K�K���K K K ����KDK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KhK�K�K���K K K ����KeK�K�K���K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KeK�K�K���K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KeK�K�K���K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KvK�K�K���K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KvK�K�K���K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KvK�K�K���K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KcK�K�K���K K K ����KeK�K�K���K K K ����KgK�K�K���K K K ����KlK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KgK�K�K���K K K ����KlK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KhK�K�K���K K K ����KeK�K�K���K K K ����KgK�K�K���K K K ����KlK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KkK�K�K���K K K ����KlK�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����KbK�K�K���K K K ����KlK�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KlK�K�K���K K K ����KeK�K�K���K K K ����KsK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KmK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K1K�K�K���K K K ����K1K�K�K���K K K ����KiK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K1K�K�K���K K K ����K5K�K�K���K K K ����KaK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K1K�K�K���K K K ����K5K�K�K���K K K ����KmK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KfK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KcK�K�K���K K K ����KuK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KfK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����KBK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KcK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KmK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KcK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KpK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KcK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����KcK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KcK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e��bub�nextSeed�M7Bub�textWall��Cracked stone wall
��	textSpace��Dusty stone floor
��djikstra_Player_Away�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�h�     G�i      G�iP     G�i�     NNNNNNNNNNNNNNNNNG�k`     G�k�     G�k�     G�k�     G�l      G�lP     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK G�n      G�m�     G�m�     G�mp     G�m@     G�m     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�h�     G�h�     G�i      G�iP     NNNNNNNNNNNNNNNNNG�k0     G�k`     G�k�     G�k�     G�k�     G�l      NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�n      G�m�     G�m�     G�mp     G�m@     G�m     G�l�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�h0     G�h`     G�h�     G�h�     G�h�     G�i      NNNNNNNNNNNNNNNNNG�k      G�k0     G�k`     G�k�     G�k�     G�k�     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�m�     G�m�     G�mp     G�m@     G�m     G�l�     G�l�     G�l�     G�lP     G�l      G�k�     G�k�     G�k�     G�k`     G�k0     G�k      NNNNNNNNNNNNNNNNNNNG�i      G�h�     G�h�     G�h�     G�h`     G�h0     G�h      G�h0     G�h`     G�h�     G�h�     G�h�     NNNNNNNNNNNNNNNNNG�j�     G�k      G�k0     G�k`     G�k�     G�k�     G�k�     G�l      G�lP     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�n      G�m�     G�m�     G�mp     G�m@     G�m     G�l�     NNNNNNNNG�j�     NNNNNNNNNNNNNNNNNNNG�iP     NNNNNG�g�     G�h      G�h0     G�h`     G�h�     G�h�     NNNNNNNNNNNNNNNNNG�j�     G�j�     G�k      G�k0     G�k`     G�k�     G�k�     G�k�     G�l      NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK G�n      G�m�     G�m�     G�mp     G�m@     G�m     NNNNNNNNG�j�     NNNNNNNNNNNNNNNNNNNG�i�     NNNNNG�g�     G�g�     G�h      G�h0     G�h`     G�h�     G�h�     G�h�     G�i      G�iP     G�i�     G�i�     G�i�     G�j     G�j@     G�jp     NNNNNNNG�jp     G�j�     G�j�     G�k      G�k0     G�k`     G�k�     G�k�     G�k�     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�n      G�m�     G�m�     G�m�     G�m�     G�mp     G�m@     NNNNNNNNG�jp     NNNNG�i�     G�iP     G�i      G�h�     G�i      G�iP     NNNNNNNNNG�i�     NNNNNG�gp     NNNNNNNNNNNNNNG�j�     G�j�     G�k      G�k0     G�k      G�j�     G�j�     G�jp     G�j@     G�jp     G�j�     G�j�     G�k      G�k0     G�k`     G�k�     G�k�     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�m�     G�m�     G�mp     G�m�     G�m�     G�m�     G�mp     NNNNNNNNG�j@     G�j     G�i�     G�i�     G�i�     G�iP     G�i      G�h�     G�h�     G�h�     G�i      G�iP     G�i�     G�i�     G�i�     G�j     G�j@     G�jp     G�j@     G�j     G�i�     NNNNNG�g@     NNNNNNNNNNNNNNNNNNNNNNG�j     G�j@     G�jp     G�j�     G�j�     G�k      G�k0     G�k`     G�k�     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�m�     G�mp     G�m@     G�mp     G�m�     G�m�     G�m�     NNNNNNNNNNNNNG�i      G�h�     G�h�     G�h�     NNNNNNNNNNNNNNNNNG�g     NNNNNNNNNNNNNNNNNNNNNNG�i�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�mp     G�m@     G�m     G�m@     G�mp     G�m�     G�m�     NNNNNNNNNNNNNG�h�     G�h�     G�h�     G�h`     NNNNNNNNNNNNNNNNNG�f�     NNNNNNNNNNNNNNNNNNNNNNG�i�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�m@     G�m     G�l�     G�m     G�m@     G�mp     G�m�     NNNNNNNNNNNNNG�h�     G�h�     G�h`     G�h0     G�h`     G�h�     NNNNNNNNNNNNNNNG�f�     NNNNNNNNNNNNNNNNNNNNNNG�i�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�l�     NNNNNNNNNNNNNNNNNG�h�     G�h`     G�h0     G�h      G�h0     G�h`     NNNNNNNNNNNNNNNG�f�     NNNNNNNNNNNNNNNNNNNNNNG�iP     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�l�     NNNNNNNNNNNNNNNNNG�h`     G�h0     G�h      G�g�     G�h      G�h0     NNNNNNNNNNNNNNNG�fP     NNNNNNNNNNNNNNNNNNNNNNG�i      NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�lP     NNNNNNNNNNNNNNNNNG�h0     G�h      G�g�     G�g�     G�g�     G�h      NNNNNNNNNNNNNNNG�f      NNNNNNNNNNNNNNNNNNNNNNG�h�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�l      NNNNNNNNNNNNNNNNNNNNG�gp     NNNNNNNNNNNNNNNNNG�e�     G�e�     G�e�     G�e`     G�e0     G�e      G�d�     NNNNNNNNNNNNNNNNG�h�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�k�     NNNNNNNNNNNNNNNNNNNNG�g@     NNNNNNNNNNNNNNNNNNNNNNNG�d�     NNNNNNNNNNNNNNNNG�h�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�k�     NNNNNNNNNNNNNNNNNNNNG�g     NNNNNNNNNNNNNNNNNNNNNNNG�dp     NNNNNNNNNNNNNNNNG�h`     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�k�     NNNNNNNNNNNNNNNNNNNNG�f�     G�f�     NNNNNNNNNNNNNNNNNNNNNNG�d@     NNNNNNNNNNNNNNNNG�h0     G�h      G�g�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�k`     NNNNNNNNNNNNNNNNNNNNNG�f�     NNNNNNNNNNNNNNNNNNNNNNG�d     NNNNNNNNNNNNNNNNNNG�g�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�j�     G�j�     G�k      G�k0     NNNNNNNNNNNNNNNNNNNNNG�fP     NNNNNNNNNNNNNNNNNNNNNNG�c�     NNNNNNNNNNNNNNNNNNG�gp     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�jp     NNNNNNNNNNNNNNNNNNG�e`     G�e0     G�e`     G�e�     G�e�     G�e�     G�f      G�fP     G�f�     G�f�     NNNNNNNNNNNNNNNNNNNG�c�     NNNNNNNNNNNNNNNNNNG�g@     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�j@     NNNNNNNNNNNNNNNNNNG�e0     G�e      G�e0     G�e`     G�e�     G�e�     G�e�     G�f      G�fP     G�f�     G�fP     G�f      G�e�     G�e�     G�e�     G�e`     G�e0     G�e      NNNNNNNNNNNG�c�     NNNNNNNNNNNNNNNNNNG�g     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�j     NNNNNNNNNNNNNNNNNNG�e      G�d�     G�e      G�e0     G�e`     G�e�     G�e�     G�e�     G�f      G�fP     NNNNNNNG�d�     NNNNNNNNNNNG�cP     NNNNNNNNNNNNNNNNNNG�f�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�j�     G�jp     G�j@     G�j     G�i�     G�i�     G�i�     G�iP     G�i�     NNNNNNNNNNNNNNG�d�     G�d�     G�d�     NNNNG�e�     G�e�     G�f      NNNNNNNG�d�     NNNNNNNNNNNG�c      NNNNNNNNNNNNNNNNG�fP     G�f�     G�f�     G�f�     G�f�     G�f�     G�g     G�g@     G�gp     G�g�     NNNNNNNNNNNNNNNNNNNe]�(NNG�jp     G�j@     G�j     G�i�     G�i�     G�i�     G�iP     G�i      G�iP     NNNNNNNNNNNNNNG�d�     G�dp     G�d�     NNNNG�e�     G�e�     G�e�     NNNNNNNG�dp     NNNNNNNNG�b�     G�b�     G�b�     G�b�     G�c      G�cP     G�c�     G�c�     G�c�     NNNNNNNNG�e�     G�e�     G�e�     G�f      G�fP     G�f�     G�f�     G�f�     G�f�     G�f�     G�g     G�g@     G�gp     NNNNNNNNNNNNNNNNNNNe]�(NNG�j@     G�j     G�i�     G�i�     G�i�     G�iP     G�i      G�h�     G�i      NNNNNNNNG�e�     G�e`     G�e0     G�e      G�d�     G�d�     G�dp     G�d@     G�dp     NNNNG�e`     G�e�     G�e�     NNNNNNNG�d@     NNNNNNNNG�b�     G�b`     G�b�     G�b�     G�b�     G�c      G�cP     G�c�     G�c�     NNNNNNNNG�e`     NNG�fP     G�f�     G�f�     G�f�     G�fP     G�f�     G�f�     G�f�     G�g     G�g@     NNNNNNNNNNNNNNNNNNNe]�(NNG�j     G�i�     G�i�     G�i�     G�iP     G�i      G�h�     G�h�     G�h�     NNNNNNNNG�e�     NNNNNG�d@     G�d     G�d@     NNNNG�e0     G�e`     G�e�     NNNNNNNG�d     G�c�     G�c�     G�c�     G�cP     G�c      G�b�     G�b�     G�b�     G�b`     G�b0     G�b`     G�b�     G�b�     G�b�     G�c      G�cP     G�c�     NNNNNNNNG�e0     NNG�f�     G�f�     G�f�     G�fP     G�f      G�fP     G�f�     G�f�     G�f�     G�g     NNNNNNNNNNNNNNNNNNNe]�(NNG�i�     G�i�     G�i�     G�iP     G�i      G�h�     G�h�     G�h�     G�h�     NNNNNNNNG�e�     NNNNNG�d     G�c�     G�d     G�d@     G�dp     G�d�     G�d�     G�e      G�e0     G�e`     NNNNNNNNNNNNNNNNG�b0     G�b      G�b0     G�b`     G�b�     G�b�     G�b�     G�c      G�cP     NNNNNNNNG�e      NNNNG�fP     G�f      G�e�     G�f      G�fP     G�f�     G�f�     G�f�     NNNNNNNNNNNNNNNNNNNe]�(NNG�j     G�i�     G�i�     NNNNG�h`     G�h�     NNNNNNNNG�f      NNNNNG�c�     G�c�     G�c�     G�d     G�d@     G�dp     G�d�     G�d�     G�e      G�e0     NNNNNNNNNNNNNNNNG�b      G�a�     G�b      G�b0     G�b`     �      G�b�     G�b�     G�b�     G�c      NNNNNNNNG�d�     NNNNG�f      G�e�     G�e�     G�e�     G�f      G�fP     G�f�     G�f�     NNNNNNNNNNNNNNNNNNNe]�(NNG�j@     G�j     G�i�     NNNNG�h0     G�h`     NNNNNNNNG�fP     NNNNNNG�c�     NNNNNNNNNNNNNNNNNNNNNNNNG�a�     G�a�     G�a�     G�b      G�b0     G�b`     G�b�     G�b�     G�b�     NNNNNNNNG�d�     NNNNNNG�e�     NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�jp     G�j@     G�j     NNNNG�h      G�h0     NNNNNNNNG�f�     NNNNNNG�cP     NNNNNNNNNNNNNNNNNNNNNNNNG�a�     G�ap     G�a�     G�a�     G�b      G�b0     G�b`     G�b�     G�b�     G�b�     G�c      G�cP     G�c�     G�c�     G�c�     G�d     G�d@     G�dp     NNNNNNG�e`     NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�j�     G�jp     G�j@     NNNNG�g�     G�h      G�h0     G�h      G�g�     G�g�     G�gp     G�g@     G�g     G�f�     G�f�     NNNNNNG�c      NNNNNNNNNNNNNNNNNNNNNNNNNG�a@     NNNNNNNNNNNNNNNNNNNNNNG�e0     G�e      G�d�     G�d�     G�dp     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�g�     NNNNNNNNNNNNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNNG�a     NNNNNNNNNNNNNNNNNNNNNNNNNNG�d@     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�gp     NNNNNNNNNNNNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNNG�`�     G�`�     G�`�     G�`P     G�`      NNNNNNNNNNNNNNNNNNNNNNG�d     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�g@     NNNNNNNNNNNNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�_�     NNNNNNNNNNNNNNNNNNNNNNG�c�     NNNNNNNNNNNNNNNNNNNNe]�(NNNNG�f      G�fP     G�f�     G�f�     G�f�     G�g     NNNNNNNNNNNNNNNNG�b`     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�_�     NNNNNNNNNNNNNNNNNNNNNNG�c�     NNNNNNNNNNNNNNNNNNNNe]�(NNNNG�e�     NNNNNNNNNNNNNNNNNNNNNG�b0     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�_      NNNNNNNNNNNNNNNNNNNNNNG�c�     NNNNNNNNNNNNNNNNNNNNe]�(NNNNG�e�     NNNNNNNNNNNNNNNNNNNNNG�b      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�^�     NNNNNNNNNNNNNNNNNNNNG�cP     G�c�     G�cP     G�c      G�cP     NNNNNNNNNNNNNNNNNNe]�(NNNNG�e�     NNNNNNNNNNNNNNNNNNNNNG�a�     NNNNNNNNNNNNNNNNNNNNNNNG�_      G�^�     G�^`     G�^      G�]�     G�^      G�^`     G�^�     G�_      NNNNNNNNNNNNNNNNNNG�c      G�cP     G�c      G�b�     G�c      NNNNNNNNNNNNNNNNNNe]�(NNNNG�e`     NNNNNNNNNNNNNNNNNNNNNG�a�     NNNNNNNNNNNNNNNNNNNNNNNG�^�     G�^`     G�^      G�]�     G�]@     G�]�     G�^      G�^`     G�^�     NNNNNNNNNNNNNNNNNNG�b�     G�c      G�b�     G�b�     G�b�     NNNNNNNNNNNNNNNNNNe]�(NNNNG�e0     NNNNNNNNNNNNNNNNNNNNG�a�     G�ap     G�a@     G�a     G�a@     G�ap     G�a�     G�a�     G�b      NNNNNNNNNNNNNNNNG�^`     G�^      G�]�     G�]@     G�\�     G�]@     G�]�     G�^      G�^`     NNNNNNNNNNNNNNNG�b0     G�b`     G�b�     G�b�     G�b�     G�b�     G�b�     G�b�     NNNNNNNNNNNNNNNNNNe]�(NNNNG�e      NNNNNNNNNNNNNNG�b�     G�b`     G�b0     G�b      G�a�     G�a�     G�ap     G�a@     G�a     G�`�     G�a     G�a@     G�ap     G�a�     G�a�     NNNNNNNNNNNNNNNNG�^      G�]�     G�]@     G�\�     G�\�     G�\�     G�]@     G�]�     G�^      NNNNNNNNNNNNNNNG�b      G�b0     G�b`     G�b�     G�b�     G�b�     G�b`     G�b�     NNNNNNNNNNNNNNNNNNe]�(NNG�e0     G�e      G�d�     G�e      G�e0     G�e`     G�e�     G�e�     G�e�     NNNNNNNNG�b�     NNNNNG�a@     G�a     G�`�     G�`�     G�`�     G�a     G�a@     G�ap     G�a�     NNNNNNNNNNNNNNNNG�]�     G�]@     G�\�     G�\�     G�\      G�\�     G�\�     G�]@     G�]�     NNNNNNNNNG�`�     G�`�     G�a     G�a@     G�ap     G�a�     G�a�     G�b      G�b0     G�b`     G�b�     G�b`     G�b0     G�b`     NNNNNNNNNNNNNNNNNNe]�(NNG�e      G�d�     G�d�     G�d�     G�e      G�e0     G�e`     G�e�     G�e�     NNNNNNNNG�b�     NNNNNG�a     G�`�     G�`�     G�`�     G�`�     G�`�     G�a     G�a@     G�ap     NNNNNNNNNNNNNNNNG�]@     G�\�     G�\�     G�\      G�[�     G�\      G�\�     G�\�     G�]@     G�]�     G�^      G�^`     G�^�     G�_      G�_�     G�_�     G�`      G�`P     G�`�     NNNNNG�b      G�b0     G�b`     G�b�     G�b`     G�b0     G�b      G�b0     NNNNNNNNNNNNNNNNNNe]�(NNG�d�     G�d�     G�dp     G�d�     G�d�     G�e      G�e0     G�e`     G�e�     NNNNNNNNG�c      NNNNNG�`�     G�`�     G�`�     G�`P     G�`�     G�`�     G�`�     G�a     G�a@     NNNNNNNNNNNNNNNNG�\�     G�\�     G�\      G�[�     G�[`     G�[�     G�\      G�\�     G�\�     NNNNNNNNNNNNNNNG�b0     G�b`     G�b�     G�b`     G�b0     G�b      G�a�     G�b      NNNNNNNNNNNNNNNNNNe]�(NNG�d�     G�dp     G�d@     NNG�d�     G�e      G�e0     G�e`     NNNNNNNNG�cP     NNNNNG�`�     G�`�     G�`P     G�`      G�`P     G�`�     G�`�     G�`�     G�a     NNNNNNNNNNNNNNNNG�\�     G�\      G�[�     G�[`     G�[      G�[`     G�[�     G�\      G�\�     NNNNNNNNNNNNNNNNNNNNNG�a�     NNNNNNNNNNNNNNNNNNNe]�(NNG�dp     G�d@     G�d     NNG�d�     G�d�     G�e      G�e0     NNNNNNNNG�c�     NNNNNG�`�     G�`P     G�`      G�_�     G�`      G�`P     G�`�     G�`�     G�`�     NNNNNNNNNNNNNNNNG�\      G�[�     G�[`     G�[      G�Z�     G�[      G�[`     G�[�     G�\      NNNNNNNNNNNNNNNNNNNNNG�ap     NNNNNNNNNNNNNNNNNNNe]�(NNG�d@     G�d     G�c�     G�d     G�d@     G�dp     G�d�     G�d�     G�e      NNNNNNNNG�c�     NNNNNG�`P     G�`      G�_�     G�_�     G�_�     G�`      G�`P     G�`�     G�`�     NNNNNNNNNNNNNNNNG�[�     G�[`     G�[      G�Z�     G�Z@     G�Z�     G�[      G�[`     G�[�     NNNNNNNNNNNNNNNNNNNNNG�a@     NNNNNNNNNNNNNNNNNNNe]�(NNG�d     G�c�     G�c�     G�c�     G�d     G�d@     G�dp     G�d�     G�d�     NNNNNNNNG�c�     NNNNNG�`      G�_�     G�_�     G�_      G�_�     G�_�     G�`      G�`P     G�`�     NNNNNNNNNNNNNNNNNNNNG�Y�     NNNNNNNNNNNNNNNG�^`     G�^�     G�_      G�_�     G�_�     G�`      G�`P     G�`�     G�`�     G�`�     G�a     NNNNNNNNNNNNNNNNNNNe]�(NNG�c�     G�c�     G�c�     G�c�     G�c�     G�d     G�d@     G�dp     G�d�     G�d�     G�e      G�e0     G�e      G�d�     G�d�     G�dp     G�d@     G�d     NNNNNG�_�     G�_�     G�_      G�^�     G�_      G�_�     G�_�     G�`      G�`P     NNNNNNNNNNNNNNNNNNNNG�Y�     NNNNNNNNNNNNNNNG�^      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNG�cP     NNNNNNNNNNNNNNNNNNNNNNNG�^`     NNNNNNNNNNNNNNNNNNNNNNNNNG�Y      NNNNNNNNNNNNNNNG�]�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNG�c      G�b�     G�b�     G�b�     G�b`     NNNNNNNNNNNNNNNNNNNG�^      NNNNNNNNNNNNNNNNNNNNNNNNNG�X�     G�X`     G�X      G�W�     G�W@     NNNNNNNNNNNG�]@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNG�b0     NNNNNNNNNNNNNNNNNNNG�]�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�V�     NNNNNNNNNNNG�\�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNG�b      NNNNNNNNNNNNNNNNNNNG�]@     G�\�     G�\�     G�\      G�[�     NNNNNNNNNNNNNNNNNNNNNNNNNG�V�     NNNNNNNNNNNG�\�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�b�     G�b�     G�b�     G�b`     G�b0     G�b      G�a�     G�a�     G�ap     G�a@     NNNNNNNNNNNNNNNNNNNNG�[`     NNNNNNNNNNNNNNNNNNNNNNNNNG�V      NNNNNNNNNNNG�\      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�b�     G�b�     G�b`     G�b0     G�b      G�a�     G�a�     G�ap     G�a@     G�a     NNNNNNNNNNNNNNNNNNNNG�[      NNNNNNNNNNNNNNNNNNNNNNNNNG�U�     NNNNNNNNNNG�[`     G�[�     G�\      G�\�     G�\�     G�]@     G�]�     G�^      G�^`     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�b�     G�b`     G�b0     G�b      G�a�     G�a�     G�ap     G�a@     G�a     G�`�     G�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     NNNNNNNNNG�[      G�Z�     G�Z@     G�Z�     G�[      NNNNNNNNNNNNNNNNNNNNNNNNG�U`     NNNNNNNNNNG�[      G�[`     G�[�     G�\      G�\�     G�\�     G�]@     G�]�     G�^      NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�b�     G�b�     G�b`     G�b0     G�b      G�a�     G�a�     G�ap     G�a@     G�a     NNNNNNNG�^`     NNNNNNNNNG�Z�     G�Z@     G�Y�     G�Z@     G�Z�     NNNNNNNNNNNNNNNNNNG�S�     G�S      G�S�     G�S�     G�T@     G�T�     G�U      NNNNNNNNNNG�Z�     G�[      G�[`     G�[�     G�\      G�\�     G�\�     G�]@     G�]�     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�b�     G�b�     G�b�     G�b`     G�b0     G�b      NNNG�a@     NNNNNNNG�^      NNNNNNNG�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y�     G�Z@     NNNNNNNNNNNNNNNNNNG�S      G�R�     G�S      G�S�     G�S�     G�T@     G�T�     G�U      G�U`     G�U�     G�V      G�V�     G�V�     G�W@     G�W�     NNG�Z@     G�Z�     G�[      G�[`     G�[�     G�\      G�\�     G�\�     G�]@     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�c      G�b�     G�b�     G�b�     G�b`     G�b0     NNNG�ap     NNNNNNNG�]�     NNNNNNNG�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�Y�     G�Y�     NNNNNNNNNNNNNNNNNNG�R�     G�R`     G�R�     G�S      G�S�     G�S�     G�T@     NNNNNNNG�X      NNG�Y�     G�Z@     G�Z�     G�[      G�[`     G�[�     G�\      G�\�     G�\�     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�cP     G�c      G�b�     G�b�     G�b�     G�b`     NNNG�a�     NNNNNNNG�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�Y      G�Y�     NNNNNNNNNNNNNNNNNNG�R`     G�R      G�R`     G�R�     G�S      G�S�     G�S�     NNNNNNNG�X`     G�X�     G�Y      G�Y�     G�Y�     G�Z@     G�Z�     G�[      G�[`     G�[�     G�\      G�\�     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�c�     G�cP     G�c      G�b�     G�b�     G�b�     G�b`     G�b0     G�b      G�a�     NNNNNNNNNNNNNNNG�Y�     G�Y�     G�Y      G�X�     G�X`     G�X�     G�Y      NNNNNNNNNNNNNNNNNNG�R      G�Q�     G�R      G�R`     G�R�     G�S      G�S�     NNNNNNNNNNG�Y�     G�Z@     G�Z�     G�[      G�[`     G�[�     G�\      G�\�     G�\�     NNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNG�Y�     G�Y      G�X�     G�X`     G�X      G�X`     G�X�     NNNNNNNNNNNNNNNNNNG�Q�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�c      NNNNNNNNNNNNNNNNNNNNNNNNG�W�     NNNNNNNNNNNNNNNNNNNNG�Q@     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�cP     NNNNNNNNNNNNNNNNNNNNNNNNG�W@     NNNNNNNNNNNNNNNNNNNNG�P�     G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�c      NNNNNNNNNNNNNNNNNNNNNNNNG�V�     NNNNNNNNNNNNNNNNNNNNG�P�     G�P      G�P�     G�P�     G�Q@     G�Q�     G�R      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNG�V�     NNNNNNNNNNNNNNNNNNNNG�P      G�O�     G�P      G�P�     G�P�     G�Q@     G�Q�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�b0     G�b`     G�b�     G�b�     NNNNNNNNNNNNNNNNNNNNNNNNG�V      NNNNNNNNNNNNNNNNNNNNNG�N�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�b      NNNNNNNNNNNNNNNNNNNNNNNNNNNG�U�     NNNNNNNNNNNNNNNNNNNNNG�N      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�a�     NNNNNNNNNNNNNNNNNNNNNNNNNG�T�     G�U      G�U`     NNNNNNNNNNNNNNNNNNNNNG�M@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�a�     NNNNNNNNNNNNNNNNNNNNNNNNNG�T@     NNNNNNNNNNNNNNNNNNNNNNNG�L�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�ap     NNNNNNNNNNNNNNNNNNNNNNNNNG�S�     NNNNNNNNNNNNNNNNNG�G@     G�H      G�H�     G�I�     G�J@     G�K      G�K�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�a@     NNNNNNNNNNNNNNNNNNNNNG�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     NNNNNNNNNNNNNNG�F�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�a@     G�a     G�`�     G�`�     G�`�     G�`P     G�`      NNNNNNNNNNNNNNNNG�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      NNNNNNNNNG�E�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�a     G�`�     G�`�     G�`�     G�`P     G�`      G�_�     NNNNNNNNNNNNNNNNG�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     NNNNG�O�     NNNNNNNNNG�E      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`�     G�`�     G�`P     G�`      G�_�     G�_�     NNNNNNNNNNNNNNNNG�U`     G�U      NNNG�S�     G�S      G�R�     NNNNG�N�     NNNNNNNNNG�D@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      NNNNNNNNNNNNNNNNG�U�     G�U`     NNNG�S�     G�S�     G�S      NNNNG�N      NNNNNNNNG�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     NNNNNNNNNNNNNNNNG�V      G�U�     NNNG�T@     G�S�     G�S�     NNNNG�M@     NNNNNNNNG�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     NNNNNNNNNNNNNNNNNG�      G�"      G�%      G�(      G�+      G�.      G�0�     G�2      G�3�     G�5      NNNNNNNNNNNNNNNNNNNe]�(NNG�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     NNNNNNNNG�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     NNNNG�L�     NNNNNNNNG�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      NNNNNNNNNNNNNNNNNG�      G�      G�"      G�%      G�(      G�+      G�.      G�0�     G�2      G�3�     NNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`P     NNG�^�     G�^`     G�^      NNNNNNNNG�Y�     NNNNNNNG�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     NNNNG�K�     NNNNNNNNG�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�(      G�%      G�"      NNNNNNG�      G�      G�      G�"      G�%      G�(      G�+      G�.      G�0�     G�2      NNNNNNNNNNNNNNNNNNNe]�(NNG�`P     G�`      NNG�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     NNNNNNNNNNNNNNNNNNNG�K      NNNNNNNNG�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      NNNNNNNNNNG�      G�      G�      G�      G��      G�       G��      G�      G�      G�      G�      G�"      G�%      G�(      G�+      G�.      G�0�     NNNNNNNNNNNNNNNNNNNe]�(NNG�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      NNNNNNNNNNNNNNNNNNNNNNNNNNNNG�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     NNNNNNNNNNNNNNNNNG�      G�      G�      G�"      G�%      G�(      G�+      G�.      G�0�     G�2      NNNNNNNNNNNNNNNNNNNe]�(NNG�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�B      G�A@     G�@�     G�?�     G�>      NNNNNNNNNNNNNNNNNG�      G�      G�"      G�%      G�(      G�+      G�.      G�0�     G�2      G�3�     NNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�B�     G�B      G�A@     G�@�     G�?�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�C�     G�B�     G�B      G�A@     G�@�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�consumeList�]�(j_  h��Bundle_Of_Arrows���h��
Gold_Coins���h�h�e�Tiles�}�(K }�(K �Tile�jp9  ��)��}�(j�  K �Objects�]�j�  j�  �row�K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K ubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�KGaj�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�Kaj�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�Kaj�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK	}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K	ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K	ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K	ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K	ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K	ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K	ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K	ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K	ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K	ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K	ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K	ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K	ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K	ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K	ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K	ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K	ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K	ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K	ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K	ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K	ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K	ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K	ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K	ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K	ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K	ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K	ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K	ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K	ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K	ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K	ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K	ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K	ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K	ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K	ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K	ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K	ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K	ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K	ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K	ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K	ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K	ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K	ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K	ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K	ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K	ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K	ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K	ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K	ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K	ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K	ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K	ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K	ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K	ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K	ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K	ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K	ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K	ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K	ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K	ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K	ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K	ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K	ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K	ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K	ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K	ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K	ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K	ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K	ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K	ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K	ubuK
}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K
ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K
ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K
ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K
ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K
ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K
ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K
ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K
ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K
ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K
ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K
ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K
ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K
ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K
ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K
ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K
ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K
ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K
ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K
ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K
ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K
ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K
ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K
ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K
ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K
ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K
ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K
ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K
ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K
ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K
ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K
ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K
ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K
ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K
ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K
ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K
ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K
ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  �       jv9  K
ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K
ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K
ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K
ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K
ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K
ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K
ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K
ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K
ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K
ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K
ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K
ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K
ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K
ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K
ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K
ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K
ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K
ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K
ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K
ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K
ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K
ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K
ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K
ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K
ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K
ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K
ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K
ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K
ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K
ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K
ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K
ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K
ubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�Kaj�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�Kaj�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  �       ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KubuK }�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K ubuK!}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K!ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K!ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K!ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K!ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K!ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K!ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K!ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K!ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K!ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K!ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K!ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K!ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K!ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K!ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K!ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K!ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K!ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K!ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K!ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K!ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K!ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K!ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K!ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K!ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K!ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K!ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K!ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K!ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K!ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K!ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K!ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K!ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K!ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K!ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K!ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K!ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K!ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K!ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K!ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K!ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K!ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K!ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K!ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K!ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K!ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K!ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K!ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K!ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K!ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K!ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K!ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K!ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K!ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K!ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K!ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K!ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K!ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K!ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K!ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K!ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K!ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K!ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K!ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K!ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K!ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K!ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K!ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K!ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K!ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K!ubuK"}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K"ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K"ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K"ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K"ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K"ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K"ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K"ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K"ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K"ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K"ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K"ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K"ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K"ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K"ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K"ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K"ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K"ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K"ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K"ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K"ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K"ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K"ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K"ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K"ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K"ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K"ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K"ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K"ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K"ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K"ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K"ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K"ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K"ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K"ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K"ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K"ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K"ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K"ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K"ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K"ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K"ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K"ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K"ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K"ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K"ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K"ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K"ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K"ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K"ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K"ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K"ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K"ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K"ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K"ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K"ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K"ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K"ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K"ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K"ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K"ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K"ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K"ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K"ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K"ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K"ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K"ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K"ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K"ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K"ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K"ubuK#}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K#ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K#ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K#ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K#ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K#ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K#ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K#ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K#ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K#ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K#ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K#ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K#ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K#ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K#ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K#ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K#ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K#ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K#ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K#ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K#ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K#ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K#ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K#ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K#ubK6jq9  )��}�(j�  K6jt9  ]�K#aj�  j�  jv9  K#ubK7jq9  )��}�(j�  K7jt9  ]�K$aj�  j�  jv9  K#ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K#ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K#ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K#ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K#ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K#ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K#ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K#ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K#ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K#ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K#ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K#ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K#ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K#ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K#ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K#ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K#ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K#ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K#ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K#ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K#ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K#ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K#ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K#ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K#ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K#ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K#ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K#ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K#ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K#ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K#ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K#ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K#ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K#ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K#ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K#ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K#ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K#ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K#ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K#ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K#ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K#ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K#ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K#ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K#ubuK$}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K$ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K$ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K$ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K$ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K$ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K$ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K$ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K$ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K$ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K$ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K$ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K$ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K$ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K$ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K$ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K$ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K$ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K$ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K$ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K$ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K$ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K$ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K$ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K$ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K$ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K$ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K$ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K$ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K$ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K$ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K$ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K$ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K$ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K$ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K$ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K$ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K$ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K$ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K$ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K$ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K$ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K$ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K$ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K$ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K$ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K$ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K$ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K$ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K$ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K$ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K$ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K$ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K$ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K$ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K$ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K$ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K$ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K$ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K$ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K$ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K$ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K$ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K$ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K$ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K$ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K$ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K$ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K$ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K$ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K$ubuK%}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K%ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K%ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K%ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K%ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K%ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K%ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K%ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K%ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K%ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K%ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K%ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K%ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K%ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K%ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K%ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K%ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K%ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K%ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K%ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K%ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K%ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K%ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K%ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K%ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K%ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K%ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K%ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K%ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K%ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K%ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K%ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K%ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K%ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K%ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K%ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K%ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K%ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K%ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K%ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K%ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K%ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K%ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K%ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K%ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K%ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K%ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K%ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K%ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K%ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K%ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K%ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K%ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K%ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K%ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K%ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K%ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K%ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K%ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K%ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K%ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K%ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K%ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K%ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K%ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K%ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K%ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K%ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K%ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K%ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K%ubuK&}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K&ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K&ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K&ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K&ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K&ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K&ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K&ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K&ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K&ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K&ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K&ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K&ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K&ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K&ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K&ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K&ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K&ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K&ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K&ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K&ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K&ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K&ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K&ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K&ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K&ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K&ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K&ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K&ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K&ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K&ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K&ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K&ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K&ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K&ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K&ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K&ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K&ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K&ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K&ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K&ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K&ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K&ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K&ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K&ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K&ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K&ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K&ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K&ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K&ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K&ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K&ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K&ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K&ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K&ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K&ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K&ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K&ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K&ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K&ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K&ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K&ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K&ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K&ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K&ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K&ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K&ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K&ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K&ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K&ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K&ubuK'}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K'ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  �      )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K'ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K'ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K'ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K'ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K'ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K'ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K'ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K'ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K'ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K'ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K'ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K'ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K'ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K'ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K'ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K'ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K'ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K'ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K'ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K'ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K'ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K'ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K'ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K'ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K'ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K'ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K'ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K'ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K'ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K'ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K'ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K'ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K'ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K'ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K'ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K'ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K'ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K'ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K'ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K'ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K'ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K'ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K'ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K'ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K'ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K'ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K'ubKNjq9  )��}�(j�  KNjt9  ]�K�aj�  j�  jv9  K'ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K'ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K'ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K'ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K'ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K'ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K'ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K'ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K'ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K'ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K'ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K'ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K'ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K'ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K'ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K'ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K'ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K'ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K'ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K'ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K'ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K'ubuK(}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K(ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K(ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K(ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K(ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K(ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K(ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K(ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K(ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K(ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K(ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K(ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K(ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K(ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K(ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K(ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K(ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K(ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K(ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K(ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K(ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K(ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K(ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K(ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K(ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K(ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K(ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K(ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K(ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K(ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K(ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K(ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K(ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K(ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K(ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K(ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K(ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K(ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K(ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K(ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K(ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K(ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K(ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K(ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K(ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K(ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K(ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K(ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K(ubKNjq9  )��}�(j�  KNjt9  ]�K'aj�  j�  jv9  K(ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K(ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K(ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K(ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K(ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K(ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K(ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K(ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K(ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K(ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K(ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K(ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K(ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K(ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K(ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K(ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K(ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K(ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K(ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K(ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K(ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K(ubuK)}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K)ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K)ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K)ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K)ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K)ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K)ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K)ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K)ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K)ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K)ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K)ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K)ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K)ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K)ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K)ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K)ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K)ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K)ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K)ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K)ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K)ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K)ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K)ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K)ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K)ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K)ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K)ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K)ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K)ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K)ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K)ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K)ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K)ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K)ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K)ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K)ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K)ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K)ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K)ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K)ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K)ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K)ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K)ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K)ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K)ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K)ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K)ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K)ubKNjq9  )��}�(j�  KNjt9  ]�K*aj�  j�  jv9  K)ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K)ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K)ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K)ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K)ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K)ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K)ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K)ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K)ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K)ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K)ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K)ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K)ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K)ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K)ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K)ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K)ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K)ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K)ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K)ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K)ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K)ubuK*}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K*ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K*ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K*ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K*ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K*ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K*ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K*ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K*ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K*ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K*ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K*ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K*ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K*ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K*ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K*ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K*ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K*ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K*ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K*ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K*ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K*ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K*ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K*ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K*ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K*ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K*ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K*ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K*ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K*ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K*ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K*ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K*ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K*ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K*ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K*ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K*ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K*ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K*ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K*ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K*ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K*ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K*ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K*ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K*ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K*ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K*ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K*ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K*ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K*ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K*ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K*ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K*ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K*ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K*ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K*ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K*ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K*ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K*ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K*ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K*ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K*ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K*ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K*ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K*ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K*ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K*ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K*ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K*ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K*ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K*ubuK+}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K+ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K+ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K+ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K+ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K+ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K+ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K+ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K+ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K+ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K+ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K+ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K+ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K+ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K+ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K+ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K+ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K+ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K+ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K+ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K+ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K+ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K+ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K+ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K+ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K+ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K+ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K+ubK9jq9  )��}�(j�  K9jt9  ]�K,aj�  j�  jv9  K+ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K+ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K+ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K+ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K+ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K+ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K+ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K+ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K+ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K+ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K+ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K+ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K+ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K+ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K+ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K+ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K+ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K+ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K+ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K+ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K+ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K+ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K+ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K+ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K+ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K+ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K+ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K+ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K+ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K+ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K+ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K+ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K+ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K+ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K+ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K+ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K+ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K+ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K+ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K+ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K+ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K+ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K+ubuK,}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�K/aj�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�K0aj�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K,ubK
jq9  )��}�(j�  K
jt9  ]�K1aj�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K,ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K,ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K,ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K,ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K,ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K,ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K,ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K,ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K,ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K,ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K,ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K,ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K,ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K,ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K,ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K,ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K,ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K,ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K,ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K,ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K,ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K,ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K,ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K,ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K,ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K,ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K,ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K,ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K,ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K,ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K,ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K,ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K,ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K,ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K,ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K,ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K,ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K,ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K,ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K,ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K,ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K,ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K,ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K,ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K,ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K,ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K,ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K,ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K,ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K,ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K,ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K,ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K,ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K,ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K,ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K,ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K,ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K,ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K,ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K,ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K,ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K,ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K,ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K,ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K,ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K,ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K,ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K,ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K,ubuK-}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K-ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�K3aj�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K-ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K-ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K-ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K-ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K-ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K-ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K-ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K-ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K-ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K-ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K-ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K-ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K-ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K-ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K-ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K-ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K-ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K-ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K-ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K-ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K-ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K-ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K-ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K-ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K-ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K-ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K-ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K-ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K-ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K-ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K-ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K-ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K-ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K-ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K-ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K-ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K-ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K-ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K-ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K-ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K-ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K-ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K-ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K-ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K-ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K-ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K-ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K-ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K-ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K-ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K-ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K-ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K-ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K-ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K-ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K-ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K-ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K-ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K-ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K-ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K-ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K-ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K-ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K-ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K-ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K-ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K-ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K-ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K-ubuK.}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K.ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K.ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K.ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K.ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K.ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K.ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K.ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K.ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K.ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K.ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K.ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K.ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K.ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K.ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K.ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K.ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K.ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K.ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K.ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K.ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K.ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K.ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K.ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K.ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K.ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K.ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K.ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K.ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K.ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K.ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K.ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K.ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K.ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K.ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K.ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K.ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K.ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K.ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K.ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K.ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K.ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K.ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K.ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K.ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K.ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K.ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K.ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K.ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K.ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K.ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K.ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K.ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K.ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K.ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K.ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K.ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K.ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K.ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K.ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K.ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K.ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K.ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K.ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K.ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K.ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K.ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K.ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K.ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K.ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K.ubuK/}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�K8aj�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K/ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K/ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K/ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K/ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K/ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K/ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K/ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K/ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K/ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K/ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K/ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K/ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K/ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K/ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K/ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K/ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K/ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K/ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K/ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K/ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K/ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K/ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K/ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K/ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K/ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K/ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K/ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K/ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K/ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K/ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K/ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K/ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K/ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K/ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K/ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K/ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K/ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K/ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K/ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K/ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K/ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K/ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K/ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K/ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K/ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K/ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K/ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K/ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K/ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K/ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K/ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K/ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K/ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K/ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K/ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K/ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K/ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K/ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K/ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K/ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K/ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K/ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K/ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K/ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K/ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K/ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K/ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K/ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K/ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K/ubuK0}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K0ubK
jq9  )��}�(j�  K
jt9  ]�K:aj�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K0ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K0ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K0ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K0ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K0ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K0ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K0ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K0ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K0ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K0ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K0ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K0ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K0ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K0ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K0ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K0ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K0ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K0ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K0ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K0ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K0ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K0ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K0ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K0ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K0ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K0ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K0ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K0ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K0ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K0ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K0ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K0ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K0ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K0ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K0ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K0ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K0ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K0ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K0ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K0ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K0ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K0ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K0ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K0ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K0ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K0ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K0ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K0ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K0ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K0ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K0ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K0ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K0ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K0ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K0ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K0ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K0ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K0ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K0ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K0ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K0ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K0ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K0ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K0ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K0ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K0ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K0ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K0ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K0ubuK1}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K1ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�K=aj�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K1ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K1ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K1ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K1ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K1ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K1ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K1ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K1ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K1ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K1ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K1ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K1ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K1ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K1ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K1ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K1ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K1ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K1ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K1ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K1ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K1ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K1ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K1ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K1ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K1ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K1ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K1ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K1ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K1ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K1ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K1ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K1ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K1ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K1ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K1ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K1ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K1ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K1ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K1ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K1ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K1ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K1ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K1ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K1ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K1ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K1ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K1ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K1ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K1ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K1ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K1ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K1ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K1ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K1ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K1ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K1ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K1ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K1ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K1ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K1ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K1ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K1ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K1ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K1ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K1ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K1ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K1ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K1ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K1ubuK2}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K2ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K2ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K2ubK!jq9  )��}�(j�  K!jt9  ]�K>aj�  j�  jv9  K2ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K2ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K2ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K2ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K2ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K2ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K2ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K2ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K2ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K2ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K2ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K2ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K2ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K2ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K2ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K2ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K2ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K2ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K2ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K2ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K2ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K2ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K2ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K2ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K2ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K2ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K2ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K2ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K2ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K2ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K2ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K2ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K2ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K2ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K2ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K2ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K2ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K2ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K2ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K2ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K2ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K2ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K2ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K2ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K2ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K2ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K2ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K2ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K2ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K2ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K2ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K2ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K2ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K2ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K2ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K2ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K2ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K2ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K2ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K2ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K2ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K2ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K2ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K2ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K2ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K2ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K2ubuK3}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K3ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K3ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K3ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K3ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K3ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K3ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K3ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K3ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K3ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K3ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K3ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K3ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K3ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K3ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K3ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K3ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K3ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K3ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K3ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K3ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K3ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K3ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K3ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K3ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K3ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K3ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K3ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K3ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K3ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K3ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K3ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K3ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K3ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K3ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K3ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K3ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K3ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K3ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K3ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K3ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K3ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K3ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K3ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K3ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K3ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K3ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K3ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K3ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K3ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K3ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K3ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K3ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K3ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K3ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K3ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K3ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K3ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K3ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K3ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K3ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K3ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K3ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K3ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K3ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K3ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K3ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K3ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K3ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K3ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K3ubuK4}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K4ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K4ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K4ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K4ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K4ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K4ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K4ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K4ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K4ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K4ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K4ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K4ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K4ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K4ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K4ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K4ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K4ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K4ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K4ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K4ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K4ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K4ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K4ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K4ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K4ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K4ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K4ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K4ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K4ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K4ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K4ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K4ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K4ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K4ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K4ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K4ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K4ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K4ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K4ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K4ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K4ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K4ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K4ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K4ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K4ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K4ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K4ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K4ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K4ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K4ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K4ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K4ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K4ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K4ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K4ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K4ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K4ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K4ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K4ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K4ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K4ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K4ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K4ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K4ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K4ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K4ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K4ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K4ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K4ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K4ubuK5}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K5ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K5ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K5ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K5ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K5ubK#jq9  )��}�(�      j�  K#jt9  ]�j�  j�  jv9  K5ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K5ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K5ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K5ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K5ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K5ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K5ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K5ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K5ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K5ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K5ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K5ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K5ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K5ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K5ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K5ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K5ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K5ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K5ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K5ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K5ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K5ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K5ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K5ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K5ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K5ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K5ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K5ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K5ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K5ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K5ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K5ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K5ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K5ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K5ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K5ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K5ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K5ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K5ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K5ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K5ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K5ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K5ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K5ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K5ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K5ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K5ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K5ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K5ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K5ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K5ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K5ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K5ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K5ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K5ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K5ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K5ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K5ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K5ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K5ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K5ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K5ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K5ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K5ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K5ubuK6}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K6ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K6ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K6ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K6ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K6ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K6ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K6ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K6ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K6ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K6ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K6ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K6ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K6ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K6ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K6ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K6ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K6ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K6ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K6ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K6ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K6ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K6ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K6ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K6ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K6ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K6ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K6ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K6ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K6ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K6ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K6ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K6ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K6ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K6ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K6ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K6ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K6ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K6ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K6ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K6ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K6ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K6ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K6ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K6ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K6ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K6ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K6ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K6ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K6ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K6ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K6ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K6ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K6ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K6ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K6ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K6ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K6ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K6ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K6ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K6ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K6ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K6ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K6ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K6ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K6ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K6ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K6ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K6ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K6ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K6ubuK7}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K7ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K7ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K7ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K7ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K7ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K7ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K7ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K7ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K7ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K7ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K7ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K7ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K7ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K7ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K7ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K7ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K7ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K7ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K7ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K7ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K7ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K7ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K7ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K7ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K7ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K7ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K7ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K7ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K7ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K7ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K7ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K7ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K7ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K7ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K7ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K7ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K7ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K7ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K7ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K7ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K7ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K7ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K7ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K7ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K7ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K7ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K7ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K7ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K7ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K7ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K7ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K7ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K7ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K7ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K7ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K7ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K7ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K7ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K7ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K7ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K7ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K7ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K7ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K7ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K7ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K7ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K7ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K7ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K7ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K7ubuK8}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K8ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K8ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K8ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K8ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K8ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K8ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K8ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K8ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K8ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K8ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K8ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K8ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K8ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K8ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K8ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K8ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K8ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K8ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K8ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K8ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K8ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K8ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K8ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K8ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K8ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K8ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K8ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K8ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K8ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K8ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K8ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K8ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K8ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K8ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K8ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K8ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K8ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K8ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K8ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K8ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K8ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K8ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K8ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K8ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K8ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K8ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K8ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K8ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K8ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K8ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K8ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K8ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K8ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K8ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K8ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K8ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K8ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K8ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K8ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K8ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K8ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K8ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K8ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K8ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K8ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K8ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K8ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K8ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K8ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K8ubuK9}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�K?aj�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�K@aj�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K9ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K9ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K9ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K9ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K9ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K9ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K9ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K9ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K9ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K9ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K9ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K9ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K9ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K9ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K9ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K9ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K9ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K9ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K9ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K9ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K9ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K9ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K9ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K9ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K9ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K9ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K9ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K9ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K9ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K9ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K9ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K9ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K9ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K9ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K9ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K9ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K9ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K9ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K9ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K9ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K9ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K9ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K9ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K9ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K9ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K9ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K9ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K9ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K9ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K9ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K9ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K9ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K9ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K9ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K9ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K9ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K9ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K9ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K9ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K9ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K9ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K9ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K9ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K9ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K9ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K9ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K9ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K9ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K9ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K9ubuK:}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K:ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K:ubKjq9  )��}�(j�  Kjt9  ]�KCaj�  j�  jv9  K:ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K:ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K:ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K:ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K:ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K:ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K:ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K:ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K:ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K:ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K:ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K:ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K:ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K:ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K:ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K:ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K:ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K:ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K:ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K:ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K:ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K:ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K:ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K:ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K:ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K:ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K:ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K:ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K:ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K:ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K:ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K:ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K:ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K:ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K:ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K:ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K:ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K:ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K:ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K:ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K:ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K:ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K:ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K:ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K:ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K:ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K:ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K:ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K:ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K:ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K:ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K:ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K:ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K:ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K:ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K:ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K:ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K:ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K:ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K:ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K:ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K:ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K:ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K:ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K:ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K:ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K:ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K:ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K:ubuK;}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K;ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K;ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K;ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K;ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K;ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K;ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K;ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K;ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K;ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K;ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K;ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K;ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K;ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K;ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K;ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K;ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K;ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K;ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K;ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K;ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K;ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K;ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K;ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K;ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K;ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K;ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K;ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K;ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K;ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K;ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K;ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K;ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K;ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K;ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K;ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K;ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K;ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K;ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K;ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K;ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K;ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K;ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K;ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K;ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K;ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K;ubKLjq9  )��}�(j�  KLjt9  ]�KDaj�  j�  jv9  K;ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K;ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K;ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K;ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K;ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K;ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K;ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K;ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K;ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K;ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K;ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K;ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K;ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K;ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K;ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K;ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K;ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K;ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K;ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K;ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K;ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K;ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K;ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K;ubuK<}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K<ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K<ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K<ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K<ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K<ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K<ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K<ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K<ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K<ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K<ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K<ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K<ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K<ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K<ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K<ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K<ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K<ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K<ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K<ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K<ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K<ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K<ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K<ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K<ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K<ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K<ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K<ubK9jq9  )��}�(j�  K9jt9  ]�KEaj�  j�  jv9  K<ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K<ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K<ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K<ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K<ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K<ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K<ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K<ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K<ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K<ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K<ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K<ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K<ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K<ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K<ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K<ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K<ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K<ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K<ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K<ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K<ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K<ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K<ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K<ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K<ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K<ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K<ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K<ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K<ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K<ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K<ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K<ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K<ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K<ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K<ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K<ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K<ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K<ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K<ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K<ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K<ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K<ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K<ubuK=}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K=ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K=ubKjq9  )��}�(j�  Kjt9  ]�KHaj�  j�  jv9  K=ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K=ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K=ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K=ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K=ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K=ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K=ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K=ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K=ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K=ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K=ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K=ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K=ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K=ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K=ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K=ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K=ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K=ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K=ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K=ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K=ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K=ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K=ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K=ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K=ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K=ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K=ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K=ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K=ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K=ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K=ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K=ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K=ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K=ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K=ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K=ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K=ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K=ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K=ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K=ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K=ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K=ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K=ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K=ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K=ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K=ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K=ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K=ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K=ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K=ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K=ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K=ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K=ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K=ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K=ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K=ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K=ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K=ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K=ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K=ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K=ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K=ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K=ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K=ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K=ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K=ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K=ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K=ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K=ubuK>}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�KBaj�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K>ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K>ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K>ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K>ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K>ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K>ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K>ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K>ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K>ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K>ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K>ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K>ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K>ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K>ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K>ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K>ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K>ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K>ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K>ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K>ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K>ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K>ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K>ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K>ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K>ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K>ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K>ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K>ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K>ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K>ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K>ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K>ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K>ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K>ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K>ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K>ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K>ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K>ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K>ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K>ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K>ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K>ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K>ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K>ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K>ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K>ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K>ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K>ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K>ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K>ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K>ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K>ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K>ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K>ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K>ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K>ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K>ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K>ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K>ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K>ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K>ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K>ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K>ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K>ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K>ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K>ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K>ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K>ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K>ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K>ubuK?}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�K9aj�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K?ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K?ubKjq9  )��}�(j�  Kjt9  ]�KLaj�  j�  jv9  K?ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K?ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K?ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K?ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K?ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K?ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K?ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K?ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K?ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K?ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K?ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K?ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K?ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K?ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K?ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K?ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K?ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K?ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K?ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K?ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K?ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K?ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K?ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K?ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K?ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K?ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K?ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K?ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K?ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K?ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K?ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K?ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K?ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K?ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K?ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K?ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K?ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K?ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K?ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K?ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K?ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K?ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K?ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K?ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K?ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K?ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K?ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K?ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K?ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K?ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K?ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K?ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K?ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K?ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K?ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K?ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K?ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K?ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K?ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K?ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K?ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K?ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K?ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K?ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K?ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K?ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K?ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K?ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K?ubuK@}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K@ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K@ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K@ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K@ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K@ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K@ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K@ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K@ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K@ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K@ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K@ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K@ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K@ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K@ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K@ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K@ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K@ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K@ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K@ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K@ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K@ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K@ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K@ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K@ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K@ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K@ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K@ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K@ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K@ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K@ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K@ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K@ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K@ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K@ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K@ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K@ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K@ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K@ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K@ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K@ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K@ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K@ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K@ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K@ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K@ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K@ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K@ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K@ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K@ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K@ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K@ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K@ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K@ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K@ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K@ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K@ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K@ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K@ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K@ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K@ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K@ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K@ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K@ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K@ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K@ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K@ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K@ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K@ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K@ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K@ubuKA}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KAubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KAubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KAubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KAubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KAubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KAubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KAubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KAubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KAubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KAubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KAubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KAubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KAubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KAubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KAubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KAubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KAubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KAubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KAubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KAubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KAubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KAubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KAubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KAubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KAubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KAubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KAubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KAubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KAubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KAubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KAubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KAubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KAubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KAubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KAubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KAubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KAubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KAubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KAubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KAubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KAubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KAubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KAubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KAubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KAubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KAubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KAubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KAubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KAubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KAubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KAubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KAubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KAubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KAubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KAubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KAubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KAubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KAubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KAubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KAubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KAubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KAubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KAubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KAubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KAubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KAubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KAubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KAubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KAubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KAubuKB}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�K.aj�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KBubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KBubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KBubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KBubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KBubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KBubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KBubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KBubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KBubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KBubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KBubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KBubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KBubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KBubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KBubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KBubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KBubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KBubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KBubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KBubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KBubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KBubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KBubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KBubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KBubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KBubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KBubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KBubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KBubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KBubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KBubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KBubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KBubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KBubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KBubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KBubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KBubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KBubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KBubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KBubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KBubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KBubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KBubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KBubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KBubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KBubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KBubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KBubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KBubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KBubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KBubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KBubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KBubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KBubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KBubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KBubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KBubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KBubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KBubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KBubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KBubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KBubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KBubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KBubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KBubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KBubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KBubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KBubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KBubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KBubuKC}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KCubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KCubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KCubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KCubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KCubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KCubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KCubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KCubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KCubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KCubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KCubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KCubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KCubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KCubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KCubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KCubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KCubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KCubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KCubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KCubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KCubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KCubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KCubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KCubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KCubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KCubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KCubK9jq9  )��}�(j�  K9jt9  �      ]�j�  j�  jv9  KCubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KCubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KCubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KCubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KCubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KCubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KCubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KCubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KCubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KCubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KCubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KCubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KCubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KCubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KCubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KCubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KCubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KCubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KCubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KCubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KCubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KCubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KCubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KCubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KCubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KCubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KCubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KCubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KCubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KCubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KCubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KCubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KCubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KCubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KCubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KCubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KCubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KCubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KCubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KCubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KCubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KCubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KCubuKD}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KDubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KDubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KDubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KDubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KDubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KDubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KDubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KDubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KDubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KDubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KDubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KDubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KDubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KDubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KDubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KDubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KDubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KDubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KDubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KDubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KDubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KDubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KDubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KDubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KDubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KDubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KDubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KDubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KDubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KDubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KDubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KDubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KDubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KDubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KDubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KDubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KDubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KDubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KDubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KDubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KDubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KDubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KDubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KDubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KDubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KDubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KDubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KDubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KDubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KDubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KDubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KDubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KDubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KDubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KDubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KDubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KDubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KDubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KDubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KDubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KDubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KDubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KDubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KDubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KDubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KDubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KDubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KDubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KDubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KDubuKE}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�KKaj�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�KWaj�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�KPaj�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KEubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KEubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KEubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KEubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KEubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KEubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KEubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KEubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KEubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KEubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KEubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KEubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KEubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KEubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KEubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KEubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KEubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KEubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KEubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KEubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KEubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KEubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KEubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KEubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KEubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KEubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KEubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KEubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KEubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KEubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KEubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KEubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KEubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KEubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KEubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KEubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KEubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KEubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KEubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KEubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KEubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KEubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KEubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KEubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KEubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KEubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KEubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KEubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KEubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KEubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KEubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KEubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KEubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KEubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KEubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KEubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KEubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KEubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KEubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KEubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KEubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KEubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KEubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KEubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KEubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KEubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KEubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KEubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KEubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KEubuKF}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KFubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KFubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KFubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KFubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KFubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KFubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KFubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KFubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KFubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KFubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KFubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KFubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KFubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KFubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KFubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KFubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KFubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KFubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KFubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KFubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KFubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KFubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KFubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KFubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KFubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KFubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KFubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KFubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KFubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KFubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KFubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KFubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KFubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KFubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KFubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KFubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KFubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KFubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KFubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KFubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KFubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KFubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KFubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KFubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KFubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KFubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KFubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KFubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KFubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KFubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KFubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KFubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KFubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KFubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KFubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KFubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KFubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KFubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KFubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KFubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KFubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KFubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KFubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KFubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KFubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KFubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KFubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KFubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KFubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KFubuKG}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�K[aj�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KGubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KGubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KGubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KGubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KGubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KGubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KGubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KGubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KGubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KGubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KGubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KGubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KGubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KGubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KGubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KGubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KGubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KGubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KGubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KGubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KGubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KGubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KGubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KGubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KGubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KGubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KGubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KGubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KGubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KGubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KGubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KGubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KGubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KGubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KGubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KGubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KGubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KGubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KGubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KGubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KGubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KGubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KGubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KGubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KGubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KGubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KGubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KGubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KGubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KGubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KGubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KGubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KGubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KGubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KGubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KGubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KGubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KGubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KGubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KGubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KGubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KGubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KGubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KGubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KGubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KGubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KGubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KGubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KGubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KGubuKH}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KHubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KHubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KHubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KHubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KHubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KHubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KHubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KHubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KHubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KHubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KHubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KHubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KHubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KHubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KHubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KHubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KHubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KHubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KHubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KHubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KHubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KHubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KHubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KHubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KHubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KHubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KHubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KHubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KHubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KHubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KHubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KHubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KHubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KHubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KHubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KHubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KHubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KHubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KHubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KHubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KHubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KHubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KHubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KHubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KHubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KHubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KHubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KHubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KHubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KHubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KHubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KHubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KHubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KHubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KHubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KHubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KHubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KHubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KHubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KHubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KHubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KHubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KHubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KHubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KHubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KHubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KHubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KHubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KHubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KHubuKI}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KIubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KIubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KIubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KIubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KIubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KIubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KIubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KIubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KIubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KIubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KIubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KIubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KIubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KIubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KIubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KIubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KIubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KIubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KIubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KIubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KIubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KIubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KIubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KIubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KIubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KIubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KIubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KIubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KIubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KIubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KIubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KIubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KIubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KIubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KIubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KIubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KIubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KIubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KIubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KIubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KIubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KIubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KIubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KIubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KIubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KIubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KIubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KIubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KIubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KIubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KIubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KIubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KIubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KIubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KIubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KIubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KIubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KIubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KIubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KIubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KIubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KIubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KIubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KIubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KIubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KIubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KIubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KIubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KIubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KIubuKJ}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KJubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�KMaj�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KJubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KJubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KJubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KJubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KJubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KJubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KJubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KJubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KJubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KJubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KJubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KJubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KJubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KJubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KJubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KJubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KJubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KJubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KJubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KJubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KJubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KJubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KJubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KJubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KJubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KJubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KJubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KJubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KJubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KJubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KJubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KJubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KJubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KJubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KJubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KJubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KJubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KJubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KJubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KJubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KJubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KJubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KJubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KJubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KJubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KJubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KJubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KJubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KJubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KJubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KJubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KJubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KJubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KJubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KJubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KJubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KJubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KJubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KJubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KJubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KJubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KJubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KJubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KJubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KJubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KJubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KJubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KJubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KJubuKK}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�KNaj�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�KOaj�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KKubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KKubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KKubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KKubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KKubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KKubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KKubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KKubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KKubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KKubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KKubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KKubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KKubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KKubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KKubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KKubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KKubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KKubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KKubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KKubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KKubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KKubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KKubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KKubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KKubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KKubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KKubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KKubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KKubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KKubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KKubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KKubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KKubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KKubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KKubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KKubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KKubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KKubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KKubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KKubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KKubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KKubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KKubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KKubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KKubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KKubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KKubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KKubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KKubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KKubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KKubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KKubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KKubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KKubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KKubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KKubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KKubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KKubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KKubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KKubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KKubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KKubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KKubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KKubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KKubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KKubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KKubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KKubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KKubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KKubuKL}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KLubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KLubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KLubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KLubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KLubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KLubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KLubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KLubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KLubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KLubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KLubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KLubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KLubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KLubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KLubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KLubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KLubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KLubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KLubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KLubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KLubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KLubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KLubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KLubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KLubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KLubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KLubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KLubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KLubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KLubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KLubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KLubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KLubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KLubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KLubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KLubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KLubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KLubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KLubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KLubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KLubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KLubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KLubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KLubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KLubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KLubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KLubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KLubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KLubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KLubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KLubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KLubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KLubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KLubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KLubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KLubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KLubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KLubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KLubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KLubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KLubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KLubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KLubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KLubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KLubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KLubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KLubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KLubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KLubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KLubuKM}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�KQaj�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KMubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KMubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KMubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KMubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KMubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KMubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KMubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KMubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KMubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KMubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KMubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KMubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KMubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KMubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KMubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KMubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KMubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KMubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KMubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KMubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KMubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KMubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KMubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KMubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KMubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KMubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KMubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KMubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KMubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KMubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KMubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KMubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KMubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KMubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KMubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KMubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KMubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KMubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KMubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KMubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KMubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KMubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KMubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KMubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KMubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KMubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KMubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KMubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KMubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KMubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KMubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KMubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KMubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KMubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KMubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KMubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KMubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KMubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KMubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KMubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KMubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KMubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KMubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KMubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KMubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KMubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KMubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KMubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KMubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KMubuKN}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�KRaj�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�KSaj�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KNubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KNubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KNubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KNubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KNubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KNubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KNubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KNubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KNubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KNubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KNubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KNubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KNubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KNubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KNubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KNubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KNubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KNubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KNubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KNubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KNubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KNubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KNubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KNubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KNubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KNubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KNubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KNubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KNubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KNubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KNubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KNubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KNubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KNubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KNubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KNubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KNubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KNubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KNubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KNubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KNubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KNubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KNubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KNubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KNubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KNubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KNubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KNubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KNubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KNubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KNubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KNubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KNubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KNubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KNubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KNubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KNubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KNubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KNubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KNubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KNubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KNubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KNubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KNubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KNubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KNubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KNubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KNubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KNubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KNubuKO}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KOubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�KTaj�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KOubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KOubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KOubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KOubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KOubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KOubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KOubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KOubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KOubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KOubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KOubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KOubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KOubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KOubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KOubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KOubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KOubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KOubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KOubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KOubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KOubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KOubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KOubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KOubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KOubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KOubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KOubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KOubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KOubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KOubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KOubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KOubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KOubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KOubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KOubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KOubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KOubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KOubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KOubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KOubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KOubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KOubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KOubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KOubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KOubKLjq9  )��}�(j�  KLjt9  ]�KVaj�  j�  jv9  KOubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KOubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KOubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KOubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KOubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KOubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KOubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KOubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KOubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KOubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KOubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KOubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KOubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KOubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KOubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KOubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KOubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KOubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KOubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KOubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KOubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KOubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KOubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KOubuKP}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KPubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�KXaj�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�KYaj�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�KZaj�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KPubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KPubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KPubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KPubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KPubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KPubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KPubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KPubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KPubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KPubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KPubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KPubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KPubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KPubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KPubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KPubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KPubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KPubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KPubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KPubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KPubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KPubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KPubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KPubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KPubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KPubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KPubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KPubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KPubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KPubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KPubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KPubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KPubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KPubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KPubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KPubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KPubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KPubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KPubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KPubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KPubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KPubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KPubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KPubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KPubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KPubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KPubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KPubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KPubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KPubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KPubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KPubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KPubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KPubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KPubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KPubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KPubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KPubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KPubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KPubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KPubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KPubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KPubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KPubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KPubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KPubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KPubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KPubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KPubuKQ}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KQubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�K]aj�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KQubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KQubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KQubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KQubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KQubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KQubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KQubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KQubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KQubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KQubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KQubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KQubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KQubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KQubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KQubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KQubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KQubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KQubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KQubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KQubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KQubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KQubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KQubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KQubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KQubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KQubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KQubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KQubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KQubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KQubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KQubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KQubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KQubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KQubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KQubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KQubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KQubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KQubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KQubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KQubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KQubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KQubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KQubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KQubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KQubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KQubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KQubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KQubKOjq9  )��}�(j�  �      KOjt9  ]�j�  j�  jv9  KQubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KQubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KQubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KQubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KQubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KQubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KQubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KQubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KQubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KQubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KQubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KQubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KQubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KQubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KQubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KQubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KQubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KQubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KQubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KQubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KQubuKR}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KRubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�Kbaj�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�Kcaj�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�Kdaj�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KRubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KRubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KRubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KRubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KRubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KRubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KRubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KRubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KRubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KRubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KRubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KRubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KRubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KRubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KRubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KRubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KRubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KRubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KRubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KRubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KRubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KRubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KRubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KRubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KRubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KRubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KRubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KRubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KRubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KRubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KRubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KRubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KRubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KRubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KRubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KRubKCjq9  )��}�(j�  KCjt9  ]�(K�K�ej�  j�  jv9  KRubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KRubKEjq9  )��}�(j�  KEjt9  ]�KFaj�  j�  jv9  KRubKFjq9  )��}�(j�  KFjt9  ]�(K�K�K�ej�  j�  jv9  KRubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KRubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KRubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KRubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KRubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KRubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KRubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KRubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KRubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KRubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KRubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KRubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KRubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KRubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KRubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KRubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KRubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KRubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KRubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KRubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KRubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KRubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KRubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KRubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KRubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KRubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KRubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KRubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KRubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KRubuKS}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KSubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KSubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KSubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KSubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KSubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KSubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KSubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KSubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KSubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KSubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KSubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KSubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KSubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KSubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KSubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KSubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KSubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KSubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KSubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KSubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KSubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KSubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KSubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KSubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KSubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KSubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KSubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KSubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KSubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KSubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KSubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KSubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KSubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KSubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KSubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KSubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KSubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KSubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KSubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KSubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KSubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KSubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KSubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KSubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KSubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KSubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KSubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KSubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KSubKOjq9  )��}�(j�  KOjt9  ]�Khaj�  j�  jv9  KSubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KSubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KSubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KSubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KSubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KSubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KSubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KSubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KSubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KSubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KSubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KSubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KSubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KSubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KSubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KSubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KSubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KSubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KSubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KSubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KSubuKT}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KTubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KTubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KTubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KTubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KTubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KTubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KTubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KTubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KTubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KTubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KTubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KTubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KTubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KTubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KTubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KTubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KTubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KTubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KTubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KTubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KTubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KTubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KTubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KTubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KTubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KTubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KTubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KTubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KTubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KTubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KTubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KTubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KTubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KTubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KTubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KTubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KTubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KTubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KTubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KTubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KTubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KTubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KTubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KTubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KTubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KTubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KTubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KTubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KTubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KTubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KTubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KTubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KTubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KTubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KTubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KTubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KTubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KTubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KTubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KTubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KTubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KTubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KTubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KTubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KTubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KTubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KTubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KTubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KTubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KTubuKU}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KUubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KUubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KUubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KUubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KUubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KUubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KUubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KUubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KUubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KUubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KUubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KUubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KUubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KUubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KUubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KUubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KUubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KUubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KUubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KUubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KUubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KUubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KUubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KUubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KUubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KUubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KUubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KUubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KUubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KUubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KUubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KUubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KUubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KUubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KUubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KUubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KUubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KUubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KUubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KUubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KUubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KUubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KUubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KUubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KUubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KUubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KUubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KUubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KUubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KUubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KUubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KUubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KUubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KUubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KUubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KUubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KUubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KUubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KUubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KUubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KUubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KUubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KUubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KUubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KUubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KUubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KUubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KUubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KUubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KUubuKV}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KVubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KVubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KVubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KVubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KVubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KVubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KVubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KVubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KVubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KVubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KVubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KVubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KVubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KVubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KVubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KVubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KVubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KVubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KVubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KVubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KVubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KVubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KVubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KVubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KVubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KVubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KVubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KVubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KVubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KVubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KVubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KVubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KVubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KVubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KVubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KVubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KVubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KVubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KVubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KVubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KVubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KVubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KVubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KVubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KVubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KVubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KVubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KVubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KVubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KVubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KVubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KVubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KVubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KVubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KVubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KVubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KVubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KVubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KVubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KVubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KVubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KVubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KVubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KVubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KVubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KVubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KVubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KVubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KVubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KVubuKW}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KWubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KWubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KWubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KWubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KWubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KWubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KWubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KWubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KWubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KWubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KWubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KWubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KWubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KWubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KWubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KWubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KWubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KWubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KWubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KWubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KWubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KWubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KWubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KWubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KWubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KWubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KWubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KWubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KWubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KWubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KWubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KWubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KWubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KWubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KWubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KWubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KWubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KWubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KWubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KWubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KWubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KWubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KWubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KWubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KWubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KWubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KWubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KWubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KWubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KWubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KWubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KWubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KWubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KWubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KWubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KWubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KWubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KWubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KWubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KWubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KWubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KWubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KWubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KWubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KWubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KWubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KWubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KWubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KWubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KWubuKX}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KXubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KXubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KXubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KXubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KXubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KXubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KXubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KXubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KXubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KXubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KXubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KXubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KXubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KXubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KXubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KXubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KXubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KXubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KXubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KXubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KXubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KXubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KXubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KXubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KXubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KXubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KXubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KXubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KXubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KXubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KXubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KXubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KXubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KXubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KXubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KXubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KXubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KXubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KXubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KXubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KXubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KXubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KXubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KXubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KXubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KXubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KXubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KXubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KXubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KXubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KXubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KXubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KXubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KXubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KXubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KXubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KXubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KXubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KXubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KXubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KXubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KXubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KXubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KXubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KXubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KXubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KXubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KXubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KXubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KXubuKY}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KYubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KYubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KYubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KYubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KYubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KYubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KYubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KYubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KYubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KYubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KYubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KYubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KYubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KYubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KYubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KYubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KYubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KYubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KYubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KYubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KYubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KYubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KYubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KYubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KYubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KYubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KYubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KYubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KYubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KYubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KYubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KYubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KYubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KYubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KYubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KYubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KYubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KYubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KYubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KYubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KYubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KYubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KYubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KYubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KYubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KYubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KYubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KYubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KYubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KYubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KYubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KYubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KYubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KYubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KYubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KYubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KYubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KYubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KYubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KYubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KYubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KYubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KYubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KYubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KYubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KYubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KYubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KYubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KYubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KYubuKZ}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KZubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KZubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KZubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KZubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KZubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KZubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KZubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KZubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KZubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KZubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KZubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KZubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KZubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KZubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KZubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KZubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KZubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KZubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KZubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KZubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KZubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KZubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KZubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KZubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KZubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KZubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KZubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KZubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KZubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KZubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KZubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KZubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KZubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KZubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KZubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KZubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KZubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KZubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KZubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KZubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KZubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KZubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KZubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KZubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KZubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KZubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KZubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KZubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KZubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KZubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KZubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KZubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KZubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KZubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KZubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KZubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KZubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KZubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KZubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KZubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KZubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KZubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KZubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KZubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KZubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KZubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KZubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KZubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KZubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KZubuK[}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K[ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K[ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K[ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K[ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K[ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K[ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K[ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K[ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K[ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K[ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K[ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K[ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K[ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K[ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K[ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K[ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K[ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K[ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K[ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K[ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K[ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K[ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K[ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K[ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K[ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K[ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K[ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K[ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K[ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K[ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K[ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K[ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K[ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K[ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K[ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K[ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K[ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K[ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K[ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K[ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K[ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K[ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K[ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K[ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K[ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K[ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K[ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K[ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K[ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K[ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K[ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K[ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K[ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K[ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K[ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K[ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K[ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K[ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K[ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K[ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K[ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K[ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K[ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K[ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K[ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K[ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K[ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K[ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K[ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K[ubuK\}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K\ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K\ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K\ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K\ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K\ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K\ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K\ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K\ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K\ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K\ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K\ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K\ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K\ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K\ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K\ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K\ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K\ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K\ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K\ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K\ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K\ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K\ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K\ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K\ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K\ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K\ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K\ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K\ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K\ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K\ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K\ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K\ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K\ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K\ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K\ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K\ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K\ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K\ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K\ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K\ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K\ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K\ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K\ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K\ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K\ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K\ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K\ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K\ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K\ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K\ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K\ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K\ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K\ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K\ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K\ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K\ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K\ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K\ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K\ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K\ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K\ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K\ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K\ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K\ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K\ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K\ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K\ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K\ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K\ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K\ubuK]}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K]ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K]ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K]ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K]ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K]ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K]ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K]ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K]ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K]ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K]ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K]ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K]ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K]ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K]ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K]ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K]ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K]ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K]ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K]ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K]ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K]ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K]ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K]ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K]ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K]ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K]ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K]ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K]ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K]ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K]ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K]ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K]ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K]ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K]ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K]ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K]ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K]ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K]ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K]ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K]ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K]ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K]ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K]ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K]ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K]ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K]ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K]ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K]ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K]ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K]ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K]ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K]ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K]ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K]ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K]ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K]ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K]ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K]ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K]ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K]ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K]ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K]ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K]ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K]ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K]ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K]ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K]ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K]ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K]ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K]ubuK^}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K^ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K^ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K^ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K^ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K^ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K^ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K^ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K^ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K^ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K^ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K^ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K^ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K^ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K^ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K^ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K^ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K^ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K^ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K^ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K^ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K^ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K^ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K^ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K^ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K^ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K^ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K^ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K^ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K^ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K^ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K^ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K^ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K^ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K^ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K^ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K^ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K^ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K^ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K^ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K^ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K^ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K^ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K^ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K^ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K^ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K^ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K^ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K^ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K^ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K^ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K^ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K^ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K^ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K^ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K^ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K^ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K^ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K^ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K^ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K^ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K^ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K^ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K^ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K^ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K^ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K^ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K^ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K^ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K^ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K^ubuK_}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K_ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K_ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K_ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K_ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K_ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K_ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K_ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K_ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K_ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K_ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K_ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K_ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K_ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K_ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K_ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K_ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K_ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K_ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K_ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K_ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K_ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K_ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K_ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K_ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K_ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K_ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K_ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K_ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K_ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K_ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K_ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K_ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K_ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K_ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K_ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K_ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K_ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K_ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K_ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K_ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K_ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K_ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K_ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K_ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K_ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K_ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K_ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K_ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K_ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K_ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K_ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K_ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K_ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K_ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K_ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K_ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K_ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K_ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K_ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K_ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K_ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K_ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K_ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K_ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K_ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K_ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K_ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K_ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K_ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K_ubuK`}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  �      ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  K`ubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  K`ubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  K`ubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  K`ubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  K`ubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  K`ubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  K`ubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  K`ubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  K`ubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  K`ubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  K`ubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  K`ubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  K`ubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  K`ubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  K`ubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  K`ubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  K`ubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  K`ubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  K`ubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  K`ubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  K`ubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  K`ubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  K`ubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  K`ubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  K`ubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  K`ubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  K`ubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  K`ubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  K`ubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  K`ubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  K`ubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  K`ubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  K`ubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  K`ubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  K`ubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  K`ubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  K`ubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  K`ubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  K`ubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  K`ubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  K`ubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  K`ubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  K`ubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  K`ubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  K`ubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  K`ubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  K`ubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  K`ubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  K`ubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  K`ubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  K`ubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  K`ubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  K`ubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  K`ubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  K`ubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  K`ubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  K`ubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  K`ubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  K`ubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  K`ubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  K`ubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  K`ubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  K`ubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  K`ubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  K`ubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  K`ubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  K`ubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  K`ubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  K`ubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  K`ubuKa}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KaubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KaubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KaubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KaubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KaubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KaubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KaubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KaubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KaubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KaubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KaubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KaubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KaubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KaubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KaubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KaubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KaubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KaubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KaubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KaubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KaubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KaubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KaubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KaubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KaubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KaubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KaubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KaubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KaubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KaubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KaubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KaubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KaubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KaubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KaubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KaubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KaubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KaubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KaubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KaubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KaubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KaubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KaubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KaubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KaubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KaubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KaubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KaubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KaubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KaubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KaubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KaubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KaubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KaubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KaubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KaubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KaubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KaubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KaubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KaubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KaubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KaubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KaubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KaubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KaubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KaubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KaubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KaubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KaubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KaubuKb}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KbubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KbubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KbubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KbubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KbubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KbubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KbubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KbubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KbubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KbubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KbubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KbubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KbubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KbubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KbubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KbubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KbubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KbubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KbubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KbubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KbubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KbubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KbubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KbubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KbubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KbubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KbubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KbubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KbubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KbubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KbubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KbubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KbubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KbubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KbubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KbubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KbubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KbubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KbubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KbubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KbubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KbubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KbubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KbubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KbubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KbubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KbubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KbubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KbubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KbubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KbubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KbubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KbubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KbubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KbubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KbubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KbubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KbubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KbubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KbubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KbubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KbubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KbubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KbubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KbubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KbubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KbubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KbubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KbubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  KbubuKc}�(K jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubK	jq9  )��}�(j�  K	jt9  ]�j�  j�  jv9  KcubK
jq9  )��}�(j�  K
jt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubKjq9  )��}�(j�  Kjt9  ]�j�  j�  jv9  KcubK jq9  )��}�(j�  K jt9  ]�j�  j�  jv9  KcubK!jq9  )��}�(j�  K!jt9  ]�j�  j�  jv9  KcubK"jq9  )��}�(j�  K"jt9  ]�j�  j�  jv9  KcubK#jq9  )��}�(j�  K#jt9  ]�j�  j�  jv9  KcubK$jq9  )��}�(j�  K$jt9  ]�j�  j�  jv9  KcubK%jq9  )��}�(j�  K%jt9  ]�j�  j�  jv9  KcubK&jq9  )��}�(j�  K&jt9  ]�j�  j�  jv9  KcubK'jq9  )��}�(j�  K'jt9  ]�j�  j�  jv9  KcubK(jq9  )��}�(j�  K(jt9  ]�j�  j�  jv9  KcubK)jq9  )��}�(j�  K)jt9  ]�j�  j�  jv9  KcubK*jq9  )��}�(j�  K*jt9  ]�j�  j�  jv9  KcubK+jq9  )��}�(j�  K+jt9  ]�j�  j�  jv9  KcubK,jq9  )��}�(j�  K,jt9  ]�j�  j�  jv9  KcubK-jq9  )��}�(j�  K-jt9  ]�j�  j�  jv9  KcubK.jq9  )��}�(j�  K.jt9  ]�j�  j�  jv9  KcubK/jq9  )��}�(j�  K/jt9  ]�j�  j�  jv9  KcubK0jq9  )��}�(j�  K0jt9  ]�j�  j�  jv9  KcubK1jq9  )��}�(j�  K1jt9  ]�j�  j�  jv9  KcubK2jq9  )��}�(j�  K2jt9  ]�j�  j�  jv9  KcubK3jq9  )��}�(j�  K3jt9  ]�j�  j�  jv9  KcubK4jq9  )��}�(j�  K4jt9  ]�j�  j�  jv9  KcubK5jq9  )��}�(j�  K5jt9  ]�j�  j�  jv9  KcubK6jq9  )��}�(j�  K6jt9  ]�j�  j�  jv9  KcubK7jq9  )��}�(j�  K7jt9  ]�j�  j�  jv9  KcubK8jq9  )��}�(j�  K8jt9  ]�j�  j�  jv9  KcubK9jq9  )��}�(j�  K9jt9  ]�j�  j�  jv9  KcubK:jq9  )��}�(j�  K:jt9  ]�j�  j�  jv9  KcubK;jq9  )��}�(j�  K;jt9  ]�j�  j�  jv9  KcubK<jq9  )��}�(j�  K<jt9  ]�j�  j�  jv9  KcubK=jq9  )��}�(j�  K=jt9  ]�j�  j�  jv9  KcubK>jq9  )��}�(j�  K>jt9  ]�j�  j�  jv9  KcubK?jq9  )��}�(j�  K?jt9  ]�j�  j�  jv9  KcubK@jq9  )��}�(j�  K@jt9  ]�j�  j�  jv9  KcubKAjq9  )��}�(j�  KAjt9  ]�j�  j�  jv9  KcubKBjq9  )��}�(j�  KBjt9  ]�j�  j�  jv9  KcubKCjq9  )��}�(j�  KCjt9  ]�j�  j�  jv9  KcubKDjq9  )��}�(j�  KDjt9  ]�j�  j�  jv9  KcubKEjq9  )��}�(j�  KEjt9  ]�j�  j�  jv9  KcubKFjq9  )��}�(j�  KFjt9  ]�j�  j�  jv9  KcubKGjq9  )��}�(j�  KGjt9  ]�j�  j�  jv9  KcubKHjq9  )��}�(j�  KHjt9  ]�j�  j�  jv9  KcubKIjq9  )��}�(j�  KIjt9  ]�j�  j�  jv9  KcubKJjq9  )��}�(j�  KJjt9  ]�j�  j�  jv9  KcubKKjq9  )��}�(j�  KKjt9  ]�j�  j�  jv9  KcubKLjq9  )��}�(j�  KLjt9  ]�j�  j�  jv9  KcubKMjq9  )��}�(j�  KMjt9  ]�j�  j�  jv9  KcubKNjq9  )��}�(j�  KNjt9  ]�j�  j�  jv9  KcubKOjq9  )��}�(j�  KOjt9  ]�j�  j�  jv9  KcubKPjq9  )��}�(j�  KPjt9  ]�j�  j�  jv9  KcubKQjq9  )��}�(j�  KQjt9  ]�j�  j�  jv9  KcubKRjq9  )��}�(j�  KRjt9  ]�j�  j�  jv9  KcubKSjq9  )��}�(j�  KSjt9  ]�j�  j�  jv9  KcubKTjq9  )��}�(j�  KTjt9  ]�j�  j�  jv9  KcubKUjq9  )��}�(j�  KUjt9  ]�j�  j�  jv9  KcubKVjq9  )��}�(j�  KVjt9  ]�j�  j�  jv9  KcubKWjq9  )��}�(j�  KWjt9  ]�j�  j�  jv9  KcubKXjq9  )��}�(j�  KXjt9  ]�j�  j�  jv9  KcubKYjq9  )��}�(j�  KYjt9  ]�j�  j�  jv9  KcubKZjq9  )��}�(j�  KZjt9  ]�j�  j�  jv9  KcubK[jq9  )��}�(j�  K[jt9  ]�j�  j�  jv9  KcubK\jq9  )��}�(j�  K\jt9  ]�j�  j�  jv9  KcubK]jq9  )��}�(j�  K]jt9  ]�j�  j�  jv9  KcubK^jq9  )��}�(j�  K^jt9  ]�j�  j�  jv9  KcubK_jq9  )��}�(j�  K_jt9  ]�j�  j�  jv9  KcubK`jq9  )��}�(j�  K`jt9  ]�j�  j�  jv9  KcubKajq9  )��}�(j�  Kajt9  ]�j�  j�  jv9  KcubKbjq9  )��}�(j�  Kbjt9  ]�j�  j�  jv9  KcubKcjq9  )��}�(j�  Kcjt9  ]�j�  j�  jv9  Kcubuu�stairsUp�]�(K<K9e�SeenMap�]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKK K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKK K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K KKKK K KKKKKKKKK K K K K K K KKKK K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKK K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKK K K KKKK K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKK K K KKK K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K KKK K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K KKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K KKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKKKKK K K K K K K K K K K K K K K K K K KKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKKKKK K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKKKKK K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K KK K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKK K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKK K K K K K K K K K KKK K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKK K K K K K K K K K KKK K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K K K K K K K KKKKKKKKKKKKK K K K K KKKK K K K K K KKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K KKKKKKKKKKKK K KKKKKK K K K K KKKK K K K K K KKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K KKKKKKKKKKKK K KKKKKK K K K K KKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKK K K K K K KK K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K KKKK K K KKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K KKKK K K KKKKKKKKKKKKK K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKK K KKKKK K K K K K KKKK K K KKKKKKKKKKKKK K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKK K KKKKKKKKKKKKKK K K K KKKK K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K KKKKKK K KKKKKKKKKKKKKK K K K KKKK K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K KKKKKK K KKKKKKKKKKKKKK K K K KKKK K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K KKK K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K KKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K ee�djikstra_Player�j9  �master_Changed_Tiles�]�(]�(KCKe]�(KBKe]�(K>Ke]�(K?Ke]�(K?Ke]�(K>Ke]�(KQKDe]�(KQKFe]�(KQKDe]�(KQKFe]�(KQKDe]�(KQKFe]�(KQKDe]�(KQKFe]�(KQKDe]�(KQKFe]�(KQKDe]�(KQKFe]�(KQKDe]�(KRKFe]�(KQKGe]�(KQKHe]�(KPKIe]�(KPKJe]�(KOKKe]�(KOKLe]�(KNKMe]�(KRKDe]�(KQKCe]�(KRKFe]�(KQKGe]�(KQKHe]�(KPKIe]�(KPKJe]�(KPKKe]�(KOKLe]�(KOKMe]�(KRKDe]�(KQKCe]�(KRKFe]�(KQKGe]�(KQKHe]�(KQKIe]�(KPKJe]�(KPKKe]�(KPKLe]�(KOKMe]�(KRKDe]�(KQKCe]�(KRKFe]�(KRKGe]�(KQKHe]�(KQKIe]�(KQKJe]�(KQKKe]�(KPKLe]�(KPKMe]�(KRKDe]�(KRKCe]�(KQKBe]�(KRKFe]�(KRKGe]�(KRKHe]�(KQKIe]�(KQKJe]�(KQKKe]�(KQKLe]�(KQKMe]�(KRKDe]�(KRKCe]�(KRKBe]�(KRKAe]�(KRK@e]�(KQK?e]�(KQK>e]�(KQK=e]�(KRKFe]�(KRKGe]�(KRKHe]�(KRKIe]�(KRKJe]�(KRKKe]�(KQKLe]�(KQKMe]�(KRKDe]�(KRKCe]�(KRKBe]�(KRKAe]�(KRK@e]�(KRK?e]�(KRKFe]�(KRKGe]�(KRKHe]�(KRKIe]�(KRKJe]�(KRKKe]�(KRKLe]�(KRKMe]�(KRKDe]�(KRKCe]�(KRKBe]�(KRKAe]�(KRK@e]�(KSK?e]�(KRKFe]�(KRKGe]�(KRKHe]�(KRKIe]�(KRKJe]�(KRKKe]�(KSKLe]�(KSKMe]�(KRKDe]�(KRKCe]�(KSKBe]�(KRKFe]�(KRKGe]�(KRKHe]�(KSKIe]�(KSKJe]�(KSKKe]�(KSKLe]�(KSKMe]�(KRKDe]�(KSKCe]�(KRKFe]�(KRKGe]�(KSKHe]�(KSKIe]�(KSKJe]�(KSKKe]�(KTKLe]�(KTKMe]�(KRKDe]�(KSKCe]�(KRKFe]�(KSKGe]�(KSKHe]�(KSKIe]�(KTKJe]�(KTKKe]�(KTKLe]�(KUKMe]�(KRKDe]�(KSKCe]�(KRKFe]�(KSKGe]�(KSKHe]�(KTKIe]�(KTKJe]�(KTKKe]�(KUKLe]�(KSKDe]�(KRKFe]�(KSKGe]�(KSKHe]�(KTKIe]�(KTKJe]�(KUKKe]�(KSKDe]�(KSKFe]�(KSKDe]�(KSKFe]�(KSKDe]�(KSKFe]�(KSKDe]�(KSKFe]�(KSKDe]�(KSKFe]�(KSKDe]�(KSKFe]�(KQKDe]�(KSKDe]�(KQKDe]�(KSKDe]�(KQKDe]�(KSKDe]�(KQKDe]�(KSKDe]�(KQKDe]�(KSKDe]�(KQKDe]�(KSKDe]�(KQKDe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKFe]�(KSKEe]�(KQKFe]�(KSKFe]�(KQKFe]�(KSKFe]�(KQKFe]�(KSKFe]�(KQKFe]�(KSKFe]�(KQKFe]�(KSKFe]�(KQKFe]�(KSKFeej�  j�  �SeesMap�]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K ee�CollisionMap�]�(]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K KKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K KKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKK KKKKKKKKKKKKKKKKKKKK KKKKKK K K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKK KKKKKKKKKKKKKKKKKKKK KKKKKK K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKK KKKKK K K K K K KKKKKKKKKK KKKKKK KKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K KKKKKK KKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKKKKKKK K K K KKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKKKKKKK K K K KKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKK K K KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KK�       KKKKK KKKKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K KKKKKKKKKKKK KKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKK KKKKKKKKKKKK KKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKKKKKKKK K K KKKKK K K KKKKKKKK KKKKKKKKKKKK KKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKKKKKKKK K K KKKKK K K KKKKKKKK KKKKKKKKK K K K K K K K K KKKKKKKKK K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK K K K K K K K K KKKKK K K KKKKKKKK KKKKKKKKK K K K K K K K K KKKKKKKKK KKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K KKKKK K K KKKKKKKK K K K K K K K K K K K K K K K K K KKKKKKKKK KKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKK KKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K KKKKK K KKKKKKKKK KKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKK KKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K KKKKK K KKKKKKKKK KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKK KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K KKKKK K KKKKKKKKK KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K KKKKK K K K K K K K K K K KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K K KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKK K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKe]�(KKK K K KKK K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKe]�(KKK K K KKK K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKK K K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K KKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKK KKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKK KKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K KKKKKKKK KKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKK KKKKKKKK KKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K KKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKK KKKKKKKK KKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKK KKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKK KKKKKKKK K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKK K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK K K K KKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK KKKKKKKKKKKKKKKKKKKKKKKKKK K K KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK KKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K K K K K KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K KKKKK KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKK K KKKK K K KKKKK KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKK K KKKK K K KKKKK KKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKK K KKKK K K KKKKK KKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K KKKKK KKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K KKK K K KKKKKKKKK KKKKKKKK K K K K K K K KKKKK KKKKKKKKK K K K K K K K K K K K K K K K K K K KKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K KKK K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKK KKKKKKKKK K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKee�itemList�]�(j_  jj9  jl9  h�h�h0�Staff���j  h0�Buckler���hshlhHh�hch�h�hxh[hShQ�Iron_Breastplate���hghh�ehWj�  �djikstra_Player_Adj�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNKOKPKQNNNNNNNNNNNNNNNNNK[K\K]K^K_K`NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKpKoKnKmKlKkKjNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKMKNKOKPNNNNNNNNNNNNNNNNNKZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKoKnKmKlKkKjKiNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKJKKKLKMKNKONNNNNNNNNNNNNNNNNKYKZK[K\K]K^NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKnKmKlKkKjKiKhKgKfKeKdKcKbKaK`K_NNNNNNNNNNNNNNNNNNNKOKNKMKLKKKJKIKJKKKLKMKNNNNNNNNNNNNNNNNNNKXKYKZK[K\K]K^K_K`NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKoKnKmKlKkKjKiNNNNNNNNK^NNNNNNNNNNNNNNNNNNNKPNNNNNKHKIKJKKKLKMNNNNNNNNNNNNNNNNNKWKXKYKZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKpKoKnKmKlKkKjNNNNNNNNK]NNNNNNNNNNNNNNNNNNNKQNNNNNKGKHKIKJKKKLKMKNKOKPKQKRKSKTKUKVNNNNNNNKVKWKXKYKZK[K\K]K^NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKqKpKoKnKmKlKkNNNNNNNNK\NNNNKWKVKUKTKUKVNNNNNNNNNKRNNNNNKFNNNNNNNNNNNNNNKWKXKYKZKYKXKWKVKUKVKWKXKYKZK[K\K]NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKrKqKpKoKnKmKlNNNNNNNNK[KZKYKXKWKVKUKTKSKTKUKVKWKXKYKXKWKVKUKTKSNNNNNKENNNNNNNNNNNNNNNNNNNNNNKTKUKVKWKXKYKZK[K\NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKsKrKqKpKoKnKmNNNNNNNNNNNNNKUKTKSKRNNNNNNNNNNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNNNKSNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKtKsKrKqKpKoKnNNNNNNNNNNNNNKTKSKRKQNNNNNNNNNNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNNNKRNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKuKtKsKrKqKpKoNNNNNNNNNNNNNKSKRKQKPKQKRNNNNNNNNNNNNNNNKBNNNNNNNNNNNNNNNNNNNNNNKQNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKtNNNNNNNNNNNNNNNNNKRKQKPKOKPKQNNNNNNNNNNNNNNNKANNNNNNNNNNNNNNNNNNNNNNKPNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKuNNNNNNNNNNNNNNNNNKQKPKOKNKOKPNNNNNNNNNNNNNNNK@NNNNNNNNNNNNNNNNNNNNNNKONNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKvNNNNNNNNNNNNNNNNNKPKOKNKMKNKONNNNNNNNNNNNNNNK?NNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKwNNNNNNNNNNNNNNNNNNNNKLNNNNNNNNNNNNNNNNNK>K=K<K;K:K9K8NNNNNNNNNNNNNNNNKMNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKxNNNNNNNNNNNNNNNNNNNNKKNNNNNNNNNNNNNNNNNNNNNNNK7NNNNNNNNNNNNNNNNKLNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKyNNNNNNNNNNNNNNNNNNNNKJNNNNNNNNNNNNNNNNNNNNNNNK6NNNNNNNNNNNNNNNNKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKxNNNNNNNNNNNNNNNNNNNNKIKHNNNNNNNNNNNNNNNNNNNNNNK5NNNNNNNNNNNNNNNNKJKIKHNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKwNNNNNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKsKtKuKvNNNNNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKrNNNNNNNNNNNNNNNNNNKKKJKIKHKGKFKEKDKCKBNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNKENNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKqNNNNNNNNNNNNNNNNNNKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKpNNNNNNNNNNNNNNNNNNKKKJKIKHKGKFKEKDKCKBNNNNNNNK8NNNNNNNNNNNK0NNNNNNNNNNNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqKpKoKnKmKlKkNNNNNNNNNNNNNNKLKKKJNNNNKEKDKCNNNNNNNK7NNNNNNNNNNNK/NNNNNNNNNNNNNNNNK@KAKBKCKBKCKDKEKFKGNNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpKoKnKmKlKkKjNNNNNNNNNNNNNNKMKLKKNNNNKFKEKDNNNNNNNK6NNNNNNNNK-K,K-K.K/K0K1K2K3NNNNNNNNK<K=K>K?K@KAKBKAKBKCKDKEKFNNNNNNNNNNNNNNNNNNNe]�(NNKqKpKoKnKmKlKkKjKiNNNNNNNNKTKSKRKQKPKOKNKMKLNNNNKGKFKENNNNNNNK5NNNNNNNNK,K+K,K-K.K/K0K1K2NNNNNNNNK;NNK@KAKBKAK@KAKBKCKDKENNNNNNNNNNNNNNNNNNNe]�(NNKpKoKnKmKlKkKjKiKhNNNNNNNNKUNNNNNKOKNKMNNNNKHKGKFNNNNNNNK4K3K2K1K0K/K.K-K,K+K*K+K,K-K.K/K0K1NNNNNNNNK:NNKAKBKAK@K?K@KAKBKCKDNNNNNNNNNNNNNNNNNNNe]�(NNKoKnKmKlKkKjKiKhKgNNNNNNNNKVNNNNNKPKOKNKMKLKKKJKIKHKGNNNNNNNNNNNNNNNNK*K)K*K+K,K-K.K/K0NNNNNNNNK9NNNNK@K?K>K?K@KAKBKCNNNNNNNNNNNNNNNNNNNe]�(NNKpKoKnNNNNKgKfNNNNNNNNKWNNNNNKQKPKOKNKMKLKKKJKIKHNNNNNNNNNNNNNNNNK)K(K)K*K+K,K-K.K/NNNNNNNNK8NNNNK?K>K=K>K?K@KAKBNNNNNNNNNNNNNNNNNNNe]�(NNKqKpKoNNNNKfKeNNNNNNNNKXNNNNNNKQNNNNNNNNNNNNNNNNNNNNNNNNK(K'K(K)K*K+K,K-K.NNNNNNNNK7NNNNNNK<NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpNNNNKeKdNNNNNNNNKYNNNNNNKRNNNNNNNNNNNNNNNNNNNNNNNNK'K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6NNNNNNK;NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqNNNNKdKcKbKaK`K_K^K]K\K[KZNNNNNNKSNNNNNNNNNNNNNNNNNNNNNNNNNK%NNNNNNNNNNNNNNNNNNNNNNK:K9K8K7K6NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKeNNNNNNNNNNNNNNNNKTNNNNNNNNNNNNNNNNNNNNNNNNNK$NNNNNNNNNNNNNNNNNNNNNNNNNNK5NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKfNNNNNNNNNNNNNNNNKUNNNNNNNNNNNNNNNNNNNNNNNNNK#K"K!K KNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKgNNNNNNNNNNNNNNNNKVNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNe]�(NNNNKmKlKkKjKiKhNNNNNNNNNNNNNNNNKWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNe]�(NNNNKnNNNNNNNNNNNNNNNNNNNNNKXNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNe]�(NNNNKoNNNNNNNNNNNNNNNNNNNNNKYNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNK0K1K0K/K0NNNNNNNNNNNNNNNNNNe]�(NNNNKpNNNNNNNNNNNNNNNNNNNNNKZNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNK/K0K/K.K/NNNNNNNNNNNNNNNNNNe]�(NNNNKqNNNNNNNNNNNNNNNNNNNNNK[NNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNK.K/K.K-K.NNNNNNNNNNNNNNNNNNe]�(NNNNKrNNNNNNNNNNNNNNNNNNNNK]K\K]K^K_K`KaKbKcNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNK*K+K,K-K.K-K,K-NNNNNNNNNNNNNNNNNNe]�(NNNNKsNNNNNNNNNNNNNNKdKcKbKaK`K_K^K]K^K_K`KaKbKcKdNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNK)K*K+K,K-K,K+K,NNNNNNNNNNNNNNNNNNe]�(NNKvKuKtKuKvKwKxKyKzNNNNNNNNKeNNNNNK_K^K_K`KaKbKcKdKeNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNK"K#K$K%K&K'K(K)K*K+K,K+K*K+NNNNNNNNNNNNNNNNNNe]�(NNKwKvKuKvKwKxKyKzK{NNNNNNNNKfNNNNNK`K_K`K_K`KaKbKcKdNNNNNNNNNNNNNNNNKKKKKKKKKKKKKKKKKK K!NNNNNK)K*K+K,K+K*K)K*NNNNNNNNNNNNNNNNNNe]�(NNKvKuKtKuKvKwKxKyKzNNNNNNNNKgNNNNNKaK`K_K^K_K`KaKbKcNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNK*K+K,K+K*K)K(K)NNNNNNNNNNNNNNNNNNe]�(NNKuKtKsNNKvKwKxKyNNNNNNNNKhNNNNNK`K_K^K]K^K_K`KaKbNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNK'NNNNNNNNNNNNNNNNNNNe]�(NNKtKsKrNNKuKvKwKxNNNNNNNNKiNNNNNK_K^K]K\K]K^K_K`KaNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNK&NNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqKrKsKtKuKvKwNNNNNNNNKjNNNNNK^K]K\K[K\K]K^K_K`NNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNK%NNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpKqKrKsKtKuKvNNNNNNNNKkNNNNNK]K\K[KZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNKKKKKKK K!K"K#K$NNNNNNNNNNNNNNNNNNNe]�(NNKqKpKoKpKqKrKsKtKuKtKsKrKqKpKoKnKmKlNNNNNK\K[KZKYKZK[K\K]K^NNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKnNNNNNNNNNNNNNNNNNNNNNNNKXNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKmKlKkKjKiNNNNNNNNNNNNNNNNNNNKWNNNNNNNNNNNNNNNNNNNNNNNNNKK
K	KKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKhNNNNNNNNNNNNNNNNNNNKVNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKgNNNNNNNNNNNNNNNNNNNKUKTKSKRKQNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKlKkKjKiKhKgKfKeKdKcNNNNNNNNNNNNNNNNNNNNKPNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKkKjKiKhKgKfKeKdKcKbNNNNNNNNNNNNNNNNNNNNKONNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKjKiKhKgKfKeKdKcKbKaK`K_K^K]K\K[KZKYNNNNNNNNNKOKNKMKNKONNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKkKjKiKhKgKfKeKdKcKbNNNNNNNKXNNNNNNNNNKNKMKLKMKNNNNNNNNNNNNNNNNNNNKKKKKK KNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKlKkKjKiKhKgNNNKcNNNNNNNKWNNNNNNNKOKNKMKLKKKLKMNNNNNNNNNNNNNNNNNNKKKKK KK KKKKKKKKNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKmKlKkKjKiKhNNNKdNNNNNNNKVNNNNNNNKNKMKLKKKJKKKLNNNNNNNNNNNNNNNNNNKKKKKK KNNNNNNNK	NNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKnKmKlKkKjKiNNNKeNNNNNNNKUKTKSKRKQKPKOKNKMKLKKKJKIKJKKNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNK
KKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKoKnKmKlKkKjKiKhKgKfNNNNNNNNNNNNNNNKLKKKJKIKHKIKJNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKlNNNNNNNNNNNNNNNNNNNNKKKJKIKHKGKHKINNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKmNNNNNNNNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNK	KKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKnNNNNNNNNNNNNNNNNNNNNNNNNKENNNNNNNNNNNNNNNNNNNNK
K	KKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKmNNNNNNNNNNNNNNNNNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNKK
K	KKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKlNNNNNNNNNNNNNNNNNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNKKK
K	KKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKhKiKjKkNNNNNNNNNNNNNNNNNNNNNNNNKBNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKgNNNNNNNNNNNNNNNNNNNNNNNNNNNKANNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKfNNNNNNNNNNNNNNNNNNNNNNNNNK>K?K@NNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKeNNNNNNNNNNNNNNNNNNNNNNNNNK=NNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKdNNNNNNNNNNNNNNNNNNNNNNNNNK<NNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKcNNNNNNNNNNNNNNNNNNNNNK?K>K=K<K;K:K9K8NNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKcKbKaK`K_K^K]NNNNNNNNNNNNNNNNK>K=K<K;K:K9K8K7K6K5K4K3K2NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKbKaK`K_K^K]K\NNNNNNNNNNNNNNNNK?K>K=K<K;K:K9K8NNNNK1NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKaK`K_K^K]K\K[NNNNNNNNNNNNNNNNK@K?NNNK;K:K9NNNNK0NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK`K_K^K]K\K[KZNNNNNNNNNNNNNNNNKAK@NNNK<K;K:NNNNK/NNNNNNNNKKKKKKK K!NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK_K^K]K\K[KZKYNNNNNNNNNNNNNNNNKBKANNNK=K<K;NNNNK.NNNNNNNNKKKKKK K!K"NNNNNNNNNNNNNNNNNK:K;K<K=K>K?K@KAKBKCNNNNNNNNNNNNNNNNNNNe]�(NNK^K]K\K[KZKYKXNNNNNNNNKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NNNNK-NNNNNNNNKKKKK K!K"K#NNNNNNNNNNNNNNNNNK9K:K;K<K=K>K?K@KAKBNNNNNNNNNNNNNNNNNNNe]�(NNK_K^NNKYKXKWNNNNNNNNKLNNNNNNNKDKCKBKAK@K?K>K=NNNNK,NNNNNNNNKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/NNNNNNK8K9K:K;K<K=K>K?K@KANNNNNNNNNNNNNNNNNNNe]�(NNK^K]NNKXKWKVKUKTKSKRKQKPKOKNKMNNNNNNNNNNNNNNNNNNNK+NNNNNNNNK KK K!K"K#K$K%NNNNNNNNNNK0K1K2K3K4K5K6K7K8K9K:K;K<K=K>K?K@NNNNNNNNNNNNNNNNNNNe]�(NNK]K\K[KZKYKXKWNNNNNNNNNNNNNNNNNNNNNNNNNNNNK*K)K(K'K&K%K$K#K"K!K K!K"K#K$K%K&NNNNNNNNNNNNNNNNNK8K9K:K;K<K=K>K?K@KANNNNNNNNNNNNNNNNNNNe]�(NNK^K]K\K[KZKYKXNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK#K$K%K&K'NNNNNNNNNNNNNNNNNK9K:K;K<K=K>K?K@KAKBNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK$K%K&K'K(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK%K&K'K(K)NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej�  j�  �
stairsDown�]�(KSKOe�djikstra_Stairs_Up�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKOKPKQKRNNNNNNNNNNNNNNNNNK\K]K^K_K`KaNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKqKpKoKnKmKlKkNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNKOKPKQNNNNNNNNNNNNNNNNNK[K\K]K^K_K`NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKpKoKnKmKlKkKjNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKLKMKNKOKPNNNNNNNNNNNNNNNNNKZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKoKnKmKlKkKjKiKhKgKfKeKdKcKbKaK`NNNNNNNNNNNNNNNNNNNKPKOKNKMKLKKKJKKKLKMKNKONNNNNNNNNNNNNNNNNKYKZK[K\K]K^K_K`KaNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKpKoKnKmKlKkKjNNNNNNNNK_NNNNNNNNNNNNNNNNNNNKQNNNNNKIKJKKKLKMKNNNNNNNNNNNNNNNNNNKXKYKZK[K\K]K^K_K`NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKqKpKoKnKmKlKkNNNNNNNNK^NNNNNNNNNNNNNNNNNNNKRNNNNNKHKIKJKKKLKMKNKOKPKQKRKSKTKUKVKWNNNNNNNKWKXKYKZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKrKqKpKoKnKmKlNNNNNNNNK]NNNNKXKWKVKUKVKWNNNNNNNNNKSNNNNNKGNNNNNNNNNNNNNNKXKYKZK[KZKYKXKWKVKWKXKYKZK[K\K]K^NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKsKrKqKpKoKnKmNNNNNNNNK\K[KZKYKXKWKVKUKTKUKVKWKXKYKZKYKXKWKVKUKTNNNNNKFNNNNNNNNNNNNNNNNNNNNNNKUKVKWKXKYKZK[K\K]NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKtKsKrKqKpKoKnNNNNNNNNNNNNNKVKUKTKSNNNNNNNNNNNNNNNNNKENNNNNNNNNNNNNNNNNNNNNNKTNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKuKtKsKrKqKpKoNNNNNNNNNNNNNKUKTKSKRNNNNNNNNNNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNNNKSNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKvKuKtKsKrKqKpNNNNNNNNNNNNNKTKSKRKQKRKSNNNNNNNNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNNNKRNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKuNNNNNNNNNNNNNNNNNKSKRKQKPKQKRNNNNNNNNNNNNNNNKBNNNNNNNNNNNNNNNNNNNNNNKQNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKvNNNNNNNNNNNNNNNNNKRKQKPKOKPKQNNNNNNNNNNNNNNNKANNNNNNNNNNNNNNNNNNNNNNKPNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKwNNNNNNNNNNNNNNNNNKQKPKOKNKOKPNNNNNNNNNNNNNNNK@NNNNNNNNNNNNNNNNNNNNNNKONNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKxNNNNNNNNNNNNNNNNNNNNKMNNNNNNNNNNNNNNNNNK?K>K=K<K;K:K9NNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKyNNNNNNNNNNNNNNNNNNNNKLNNNNNNNNNNNNNNNNNNNNNNNK8NNNNNNNNNNNNNNNNKMNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKzNNNNNNNNNNNNNNNNNNNNKKNNNNNNNNNNNNNNNNNNNNNNNK7NNNNNNNNNNNNNNNNKLNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKyNNNNNNNNNNNNNNNNNNNNKJKINNNNNNNNNNNNNNNNNNNNNNK6NNNNNNNNNNNNNNNNKKKJKINNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKxNNNNNNNNNNNNNNNNNNNNNKHNNNNNNNNNNNNNNNNNNNNNNK5NNNNNNNNNNNNNNNNNNKHNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKtKuKvKwNNNNNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKsNNNNNNNNNNNNNNNNNNKLKKKJKIKHKGKFKEKDKCNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKrNNNNNNNNNNNNNNNNNNKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNKENNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKqNNNNNNNNNNNNNNNNNNKLKKKJKIKHKGKFKEKDKCNNNNNNNK9NNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKtKsKrKqKpKoKnKmKlNNNNNNNNNNNNNNKMKLKKNNNNKFKEKDNNNNNNNK8NNNNNNNNNNNK0NNNNNNNNNNNNNNNNKAKBKCKDKCKDKEKFKGKHNNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqKpKoKnKmKlKkNNNNNNNNNNNNNNKNKMKLNNNNKGKFKENNNNNNNK7NNNNNNNNK.K-K.K/K0K1K2K3K4NNNNNNNNK=K>K?K@KAKBKCKBKCKDKEKFKGNNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpKoKnKmKlKkKjNNNNNNNNKUKTKSKRKQKPKOKNKMNNNNKHKGKFNNNNNNNK6NNNNNNNNK-K,K-K.K/K0K1K2K3NNNNNNNNK<NNKAKBKCKBKAKBKCKDKEKFNNNNNNNNNNNNNNNNNNNe]�(NNKqKpKoKnKmKlKkKjKiNNNNNNNNKVNNNNNKPKOKNNNNNKIKHKGNNNNNNNK5K4K3K2K1K0K/K.K-K,K+K,K-K.K/K0K1K2NNNNNNNNK;NNKBKCKBKAK@KAKBKCKDKENNNNNNNNNNNNNNNNNNNe]�(NNKpKoKnKmKlKkKjKiKhNNNNNNNNKWNNNNNKQKPKOKNKMKLKKKJKIKHNNNNNNNNNNNNNNNNK+K*K+K,K-K.K/K0K1NNNNNNNNK:NNNNKAK@K?K@KAKBKCKDNNNNNNNNNNNNNNNNNNNe]�(NNKqKpKoNNNNKhKgNNNNNNNNKXNNNNNKRKQKPKOKNKMKLKKKJKINNNNNNNNNNNNNNNNK*K)K*K+K,K-K.K/K0NNNNNNNNK9NNNNK@K?K>K?K@KAKBKCNNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpNNNNKgKfNNNNNNNNKYNNNNNNKRNNNNNNNNNNNNNNNNNNNNNNNNK)K(K)K*K+K,K-K.K/NNNNNNNNK8NNNNNNK=NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqNNNNKfKeNNNNNNNNKZNNNNNNKSNNNNNNNNNNNNNNNNNNNNNNNNK(K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7NNNNNNK<NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKtKsKrNNNNKeKdKcKbKaK`K_K^K]K\K[NNNNNNKTNNNNNNNNNNNNNNNNNNNNNNNNNK&NNNNNNNNNNNNNNNNNNNNNNK;K:K9K8K7NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKfNNNNNNNNNNNNNNNNKUNNNNNNNNNNNNNNNNNNNNNNNNNK%NNNNNNNNNNNNNNNNNNNNNNNNNNK6NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKgNNNNNNNNNNNNNNNNKVNNNNNNNNNNNNNNNNNNNNNNNNNK$K#K"K!K NNNNNNNNNNNNNNNNNNNNNNK5NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKhNNNNNNNNNNNNNNNNKWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNNNe]�(NNNNKnKmKlKkKjKiNNNNNNNNNNNNNNNNKXNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNe]�(NNNNKoNNNNNNNNNNNNNNNNNNNNNKYNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNe]�(NNNNKpNNNNNNNNNNNNNNNNNNNNNKZNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNK1K2K1K0K1NNNNNNNNNNNNNNNNNNe]�(NNNNKqNNNNNNNNNNNNNNNNNNNNNK[NNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNK0K1K0K/K0NNNNNNNNNNNNNNNNNNe]�(NNNNKrNNNNNNNNNNNNNNNNNNNNNK\NNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNK/K0K/K.K/NNNNNNNNNNNNNNNNNNe]�(NNNNKsNNNNNNNNNNNNNNNNNNNNK^K]K^K_K`KaKbKcKdNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNK+K,K-K.K/K.K-K.NNNNNNNNNNNNNNNNNNe]�(NNNNKtNNNNNNNNNNNNNNKeKdKcKbKaK`K_K^K_K`KaKbKcKdKeNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNK*K+K,K-K.K-K,K-NNNNNNNNNNNNNNNNNNe]�(NNKwKvKuKvKwKxKyKzK{NNNNNNNNKfNNNNNK`K_K`KaKbKcKdKeKfNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNK#K$K%K&K'K(K)K*K+K,K-K,K+K,NNNNNNNNNNNNNNNNNNe]�(NNKxKwKvKwKxKyKzK{K|NNNNNNNNKgNNNNNKaK`KaK`KaKbKcKdKeNNNNNNNNNNNNNNNNKKKKKKKKKKKKKKKKK K!K"NNNNNK*K+K,K-K,K+K*K+NNNNNNNNNNNNNNNNNNe]�(NNKwKvKuKvKwKxKyKzK{NNNNNNNNKhNNNNNKbKaK`K_K`KaKbKcKdNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNK+K,K-K,K+K*K)K*NNNNNNNNNNNNNNNNNNe]�(NNKvKuKtNNKwKxKyKzNNNNNNNNKiNNNNNKaK`K_K^K_K`KaKbKcNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNK(NNNNNNNNNNNNNNNNNNNe]�(NNKuKtKsNNKvKwKxKyNNNNNNNNKjNNNNNK`K_K^K]K^K_K`KaKbNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNK'NNNNNNNNNNNNNNNNNNNe]�(NNKtKsKrKsKtKuKvKwKxNNNNNNNNKkNNNNNK_K^K]K\K]K^K_K`KaNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNK&NNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqKrKsKtKuKvKwNNNNNNNNKlNNNNNK^K]K\K[K\K]K^K_K`NNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNKKKKKK K!K"K#K$K%NNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpKqKrKsKtKuKvKuKtKsKrKqKpKoKnKmNNNNNK]K\K[KZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKoNNNNNNNNNNNNNNNNNNNNNNNKYNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKnKmKlKkKjNNNNNNNNNNNNNNNNNNNKXNNNNNNNNNNNNNNNNNNNNNNNNNKKK
K	KNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKiNNNNNNNNNNNNNNNNNNNKWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKhNNNNNNNNNNNNNNNNNNNKVKUKTKSKRNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKmKlKkKjKiKhKgKfKeKdNNNNNNNNNNNNNNNNNNNNKQNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKlKkKjKiKhKgKfKeKdKcNNNNNNNNNNNNNNNNNNNNKPNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKkKjKiKhKgKfKeKdKcKbKaK`K_K^K]K\K[KZNNNNNNNNNKPKOKNKOKPNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKlKkKjKiKhKgKfKeKdKcNNNNNNNKYNNNNNNNNNKOKNKMKNKONNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKmKlKkKjKiKhNNNKdNNNNNNNKXNNNNNNNKPKOKNKMKLKMKNNNNNNNNNNNNNNNNNNNKKKKKK KKKKKKKKK	NNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKnKmKlKkKjKiNNNKeNNNNNNNKWNNNNNNNKOKNKMKLKKKLKMNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNK
NNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKoKnKmKlKkKjNNNKfNNNNNNNKVKUKTKSKRKQKPKOKNKMKLKKKJKKKLNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNKKKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKpKoKnKmKlKkKjKiKhKgNNNNNNNNNNNNNNNKMKLKKKJKIKJKKNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKmNNNNNNNNNNNNNNNNNNNNKLKKKJKIKHKIKJNNNNNNNNNNNNNNNNNNK	KKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKnNNNNNNNNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNK
K	KKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKoNNNNNNNNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNKK
K	KKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKnNNNNNNNNNNNNNNNNNNNNNNNNKENNNNNNNNNNNNNNNNNNNNKKK
K	KKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKmNNNNNNNNNNNNNNNNNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNKKKK
K	KK	NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKiKjKkKlNNNNNNNNNNNNNNNNNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKhNNNNNNNNNNNNNNNNNNNNNNNNNNNKBNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKgNNNNNNNNNNNNNNNNNNNNNNNNNK?K@KANNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKfNNNNNNNNNNNNNNNNNNNNNNNNNK>NNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKeNNNNNNNNNNNNNNNNNNNNNNNNNK=NNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKdNNNNNNNNNNNNNNNNNNNNNK@K?K>K=K<K;K:K9NNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKdKcKbKaK`K_K^NNNNNNNNNNNNNNNNK?K>K=K<K;K:K9K8K7K6K5K4K3NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKcKbKaK`K_K^K]NNNNNNNNNNNNNNNNK@K?K>K=K<K;K:K9NNNNK2NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKbKaK`K_K^K]K\NNNNNNNNNNNNNNNNKAK@NNNK<K;K:NNNNK1NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKaK`K_K^K]K\K[NNNNNNNNNNNNNNNNKBKANNNK=K<K;NNNNK0NNNNNNNNKKKKKK K!K"NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK`K_K^K]K\K[KZNNNNNNNNNNNNNNNNKCKBNNNK>K=K<NNNNK/NNNNNNNNKKKKK K!K"K#NNNNNNNNNNNNNNNNNK;K<K=K>K?K@KAKBKCKDNNNNNNNNNNNNNNNNNNNe]�(NNK_K^K]K\K[KZKYNNNNNNNNKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=NNNNK.NNNNNNNNKKKK K!K"K#K$NNNNNNNNNNNNNNNNNK:K;K<K=K>K?K@KAKBKCNNNNNNNNNNNNNNNNNNNe]�(NNK`K_NNKZKYKXNNNNNNNNKMNNNNNNNKEKDKCKBKAK@K?K>NNNNK-NNNNNNNNK KK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0NNNNNNK9K:K;K<K=K>K?K@KAKBNNNNNNNNNNNNNNNNNNNe]�(NNK_K^NNKYKXKWKVKUKTKSKRKQKPKOKNNNNNNNNNNNNNNNNNNNNK,NNNNNNNNK!K K!K"K#K$K%K&NNNNNNNNNNK1K2K3K4K5K6K7K8K9K:K;K<K=K>K?K@KANNNNNNNNNNNNNNNNNNNe]�(NNK^K]K\K[KZKYKXNNNNNNNNNNNNNNNNNNNNNNNNNNNNK+K*K)K(K'K&K%K$K#K"K!K"K#K$K%K&K'NNNNNNNNNNNNNNNNNK9K:K;K<K=K>K?K@KAKBNNNNNNNNNNNNNNNNNNNe]�(NNK_K^K]K\K[KZKYNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK$K%K&K'K(NNNNNNNNNNNNNNNNNK:K;K<K=K>K?K@KAKBKCNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK%K&K'K(K)NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK&K'K(K)K*NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�maze�]�(]�(�#�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �.�j��  j��  �x�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �=�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  h<j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jb  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �~�j�  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jb  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  h<j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  jb  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  h<j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  �       j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �S�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j�  j�  j�  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j�  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j�  j�  j�  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  h<j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �E�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  h<j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  ee�	enemyList�]�(�Enemies.Goblins��Goblin_Stonewall���j`�  �Goblin_Lancer���j`�  �Goblin_Berserker���j`�  �Goblin_Archer���j`�  �Goblin_Knight���j`�  �Goblin_Grunt���j`�  �Goblin_Thief���e�djikstra_Stairs_Down�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK�K�K�K�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK�K�K�K�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNK�K�K�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNK�NNNNNNNNNNNNNNNNNNNK�NNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNK�NNNNNNNNNNNNNNNNNNNK�NNNNNK�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�NNNNNNNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNK�NNNNK�K�K�K�K�K�NNNNNNNNNK�NNNNNK�NNNNNNNNNNNNNNK�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNK�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�NNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNK�K�K�K�NNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNK�K�K�K�NNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNK�KK~K}K|K{KzNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNKyNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNKxNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNK�K�NNNNNNNNNNNNNNNNNNNNNNKwNNNNNNNNNNNNNNNNK�K�K�NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNKvNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�K�K�K�NNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNKuNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNK}K|K}K~KK�K�K�K�K�NNNNNNNNNNNNNNNNNNNKtNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNK|K{K|K}K~KK�K�K�K�K�K�K�KK~K}K|K{NNNNNNNNNNNKsNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNK{KzK{K|K}K~KK�K�K�NNNNNNNKzNNNNNNNNNNNKrNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNKzKyKzNNNNKK�K�NNNNNNNKyNNNNNNNNNNNKqNNNNNNNNNNNNNNNNK�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNKyKxKyNNNNK~KK�NNNNNNNKxNNNNNNNNKoKnKoKpKqKrKsKtKuNNNNNNNNK~KK�K�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK~K}K|K{KzKyKxKwKxNNNNK}K~KNNNNNNNKwNNNNNNNNKnKmKnKoKpKqKrKsKtNNNNNNNNK}NNK�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNKNNNNNKwKvKwNNNNK|K}K~NNNNNNNKvKuKtKsKrKqKpKoKnKmKlKmKnKoKpKqKrKsNNNNNNNNK|NNK�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK�NNNNNKvKuKvKwKxKyKzK{K|K}NNNNNNNNNNNNNNNNKlKkKlKmKnKoKpKqKrNNNNNNNNK{NNNNK�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK�K�NNNNNNNNK�NNNNNKuKtKuKvKwKxKyKzK{K|NNNNNNNNNNNNNNNNKkKjKkKlKmKnKoKpKqNNNNNNNNKzNNNNK�K�KK�K�K�K�K�NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK�K�NNNNNNNNK�NNNNNNKsNNNNNNNNNNNNNNNNNNNNNNNNKjKiKjKkKlKmKnKoKpNNNNNNNNKyNNNNNNK~NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK�K�NNNNNNNNK�NNNNNNKrNNNNNNNNNNNNNNNNNNNNNNNNKiKhKiKjKkKlKmKnKoKpKqKrKsKtKuKvKwKxNNNNNNK}NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK�K�K�K�K�K�K�K�K�K�K�NNNNNNKqNNNNNNNNNNNNNNNNNNNNNNNNNKgNNNNNNNNNNNNNNNNNNNNNNK|K{KzKyKxNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNKpNNNNNNNNNNNNNNNNNNNNNNNNNKfNNNNNNNNNNNNNNNNNNNNNNNNNNKwNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNKoNNNNNNNNNNNNNNNNNNNNNNNNNKeKdKcKbKaNNNNNNNNNNNNNNNNNNNNNNKvNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNKnNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK`NNNNNNNNNNNNNNNNNNNNNNKuNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNNKmNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK_NNNNNNNNNNNNNNNNNNNNNNKtNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNNKlNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK^NNNNNNNNNNNNNNNNNNNNNNKsNNNNNNNNNNNNNNNNNNNNe]�(NNNNKNNNNNNNNNNNNNNNNNNNNNKkNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK]NNNNNNNNNNNNNNNNNNNNKrKsKrKqKrNNNNNNNNNNNNNNNNNNe]�(NNNNK~NNNNNNNNNNNNNNNNNNNNNKjNNNNNNNNNNNNNNNNNNNNNNNK^K]K\K[KZK[K\K]K^NNNNNNNNNNNNNNNNNNKqKrKqKpKqNNNNNNNNNNNNNNNNNNe]�(NNNNK}NNNNNNNNNNNNNNNNNNNNNKiNNNNNNNNNNNNNNNNNNNNNNNK]K\K[KZKYKZK[K\K]NNNNNNNNNNNNNNNNNNKpKqKpKoKpNNNNNNNNNNNNNNNNNNe]�(NNNNK|NNNNNNNNNNNNNNNNNNNNKiKhKgKfKgKhKiKjKkNNNNNNNNNNNNNNNNK\K[KZKYKXKYKZK[K\NNNNNNNNNNNNNNNKlKmKnKoKpKoKnKoNNNNNNNNNNNNNNNNNNe]�(NNNNK{NNNNNNNNNNNNNNKnKmKlKkKjKiKhKgKfKeKfKgKhKiKjNNNNNNNNNNNNNNNNK[KZKYKXKWKXKYKZK[NNNNNNNNNNNNNNNKkKlKmKnKoKnKmKnNNNNNNNNNNNNNNNNNNe]�(NNK|K{KzK{K|K}K~KK�NNNNNNNNKoNNNNNKgKfKeKdKeKfKgKhKiNNNNNNNNNNNNNNNNKZKYKXKWKVKWKXKYKZNNNNNNNNNKdKeKfKgKhKiKjKkKlKmKnKmKlKmNNNNNNNNNNNNNNNNNNe]�(NNK{KzKyKzK{K|K}K~KNNNNNNNNKpNNNNNKfKeKdKcKdKeKfKgKhNNNNNNNNNNNNNNNNKYKXKWKVKUKVKWKXKYKZK[K\K]K^K_K`KaKbKcNNNNNKkKlKmKnKmKlKkKlNNNNNNNNNNNNNNNNNNe]�(NNKzKyKxKyKzK{K|K}K~NNNNNNNNKqNNNNNKeKdKcKbKcKdKeKfKgNNNNNNNNNNNNNNNNKXKWKVKUKTKUKVKWKXNNNNNNNNNNNNNNNKlKmKnKmKlKkKjKkNNNNNNNNNNNNNNNNNNe]�(NNKyKxKwNNKzK{K|K}NNNNNNNNKrNNNNNKdKcKbKaKbKcKdKeKfNNNNNNNNNNNNNNNNKWKVKUKTKSKTKUKVKWNNNNNNNNNNNNNNNNNNNNNKiNNNNNNNNNNNNNNNNNNNe]�(NNKxKwKvNNKyKzK{K|NNNNNNNNKsNNNNNKcKbKaK`KaKbKcKdKeNNNNNNNNNNNNNNNNKVKUKTKSKRKSKTKUKVNNNNNNNNNNNNNNNNNNNNNKhNNNNNNNNNNNNNNNNNNNe]�(NNKwKvKuKvKwKxKyKzK{NNNNNNNNKtNNNNNKbKaK`K_K`KaKbKcKdNNNNNNNNNNNNNNNNKUKTKSKRKQKRKSKTKUNNNNNNNNNNNNNNNNNNNNNKgNNNNNNNNNNNNNNNNNNNe]�(NNKvKuKtKuKvKwKxKyKzNNNNNNNNKuNNNNNKaK`K_K^K_K`KaKbKcNNNNNNNNNNNNNNNNNNNNKPNNNNNNNNNNNNNNNK\K]K^K_K`KaKbKcKdKeKfNNNNNNNNNNNNNNNNNNNe]�(NNKuKtKsKtKuKvKwKxKyKzK{K|K{KzKyKxKwKvNNNNNK`K_K^K]K^K_K`KaKbNNNNNNNNNNNNNNNNNNNNKONNNNNNNNNNNNNNNK[NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKrNNNNNNNNNNNNNNNNNNNNNNNK\NNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKZNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKqKpKoKnKmNNNNNNNNNNNNNNNNNNNK[NNNNNNNNNNNNNNNNNNNNNNNNNKMKLKKKJKINNNNNNNNNNNKYNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKlNNNNNNNNNNNNNNNNNNNKZNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKHNNNNNNNNNNNKXNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKkNNNNNNNNNNNNNNNNNNNKYKXKWKVKUNNNNNNNNNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNKWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKpKoKnKmKlKkKjKiKhKgNNNNNNNNNNNNNNNNNNNNKTNNNNNNNNNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNKVNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKoKnKmKlKkKjKiKhKgKfNNNNNNNNNNNNNNNNNNNNKSNNNNNNNNNNNNNNNNNNNNNNNNNKENNNNNNNNNNKTKUKVKWKXKYKZK[K\NNNNNNNNNNNNNNNNNNNNNNe]�(NNKnKmKlKkKjKiKhKgKfKeKdKcKbKaK`K_K^K]NNNNNNNNNKSKRKQKRKSNNNNNNNNNNNNNNNNNNNNNNNNKDNNNNNNNNNNKSKTKUKVKWKXKYKZK[NNNNNNNNNNNNNNNNNNNNNNe]�(NNKoKnKmKlKkKjKiKhKgKfNNNNNNNK\NNNNNNNNNKRKQKPKQKRNNNNNNNNNNNNNNNNNNK?K>K?K@KAKBKCNNNNNNNNNNKRKSKTKUKVKWKXKYKZNNNNNNNNNNNNNNNNNNNNNNe]�(NNKpKoKnKmKlKkNNNKgNNNNNNNK[NNNNNNNKSKRKQKPKOKPKQNNNNNNNNNNNNNNNNNNK>K=K>K?K@KAKBKCKDKEKFKGKHKIKJNNKQKRKSKTKUKVKWKXKYNNNNNNNNNNNNNNNNNNNNNNe]�(NNKqKpKoKnKmKlNNNKhNNNNNNNKZNNNNNNNKRKQKPKOKNKOKPNNNNNNNNNNNNNNNNNNK=K<K=K>K?K@KANNNNNNNKKNNKPKQKRKSKTKUKVKWKXNNNNNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpKoKnKmNNNKiNNNNNNNKYKXKWKVKUKTKSKRKQKPKOKNKMKNKONNNNNNNNNNNNNNNNNNK<K;K<K=K>K?K@NNNNNNNKLKMKNKOKPKQKRKSKTKUKVKWNNNNNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqKpKoKnKmKlKkKjNNNNNNNNNNNNNNNKPKOKNKMKLKMKNNNNNNNNNNNNNNNNNNNK;K:K;K<K=K>K?NNNNNNNNNNKPKQKRKSKTKUKVKWKXNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKpNNNNNNNNNNNNNNNNNNNNKOKNKMKLKKKLKMNNNNNNNNNNNNNNNNNNK:K9K:K;K<K=K>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKqNNNNNNNNNNNNNNNNNNNNNNNNKJNNNNNNNNNNNNNNNNNNNNK9K8K9K:K;K<K=NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKrNNNNNNNNNNNNNNNNNNNNNNNNKINNNNNNNNNNNNNNNNNNNNK8K7K8K9K:K;K<NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKqNNNNNNNNNNNNNNNNNNNNNNNNKHNNNNNNNNNNNNNNNNNNNNK7K6K7K8K9K:K;NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKpNNNNNNNNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNK6K5K6K7K8K9K:NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKlKmKnKoNNNNNNNNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKkNNNNNNNNNNNNNNNNNNNNNNNNNNNKENNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKjNNNNNNNNNNNNNNNNNNNNNNNNNKBKCKDNNNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKiNNNNNNNNNNNNNNNNNNNNNNNNNKANNNNNNNNNNNNNNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKhNNNNNNNNNNNNNNNNNNNNNNNNNK@NNNNNNNNNNNNNNNNNK*K+K,K-K.K/K0NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKgNNNNNNNNNNNNNNNNNNNNNKCKBKAK@K?K>K=K<NNNNNNNNNNNNNNK)NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKgKfKeKdKcKbKaNNNNNNNNNNNNNNNNKBKAK@K?K>K=K<K;K:K9K8K7K6NNNNNNNNNK(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKfKeKdKcKbKaK`NNNNNNNNNNNNNNNNKCKBKAK@K?K>K=K<NNNNK5NNNNNNNNNK'NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKeKdKcKbKaK`K_NNNNNNNNNNNNNNNNKDKCNNNK?K>K=NNNNK4NNNNNNNNNK&NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKdKcKbKaK`K_K^NNNNNNNNNNNNNNNNKEKDNNNK@K?K>NNNNK3NNNNNNNNK&K%K$K#K"K!K KNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKcKbKaK`K_K^K]NNNNNNNNNNNNNNNNKFKENNNKAK@K?NNNNK2NNNNNNNNK%K$K#K"K!K KKNNNNNNNNNNNNNNNNNKKK
K	KKKKKKNNNNNNNNNNNNNNNNNNNe]�(NNKbKaK`K_K^K]K\NNNNNNNNKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@NNNNK1NNNNNNNNK$K#K"K!K KKKNNNNNNNNNNNNNNNNNKK
K	KKKKKKKNNNNNNNNNNNNNNNNNNNe]�(NNKcKbNNK]K\K[NNNNNNNNKPNNNNNNNKHKGKFKEKDKCKBKANNNNK0NNNNNNNNK#K"K!K KKKKKKKKKKKKKKKNNNNNNK
K	KKKKKKKKNNNNNNNNNNNNNNNNNNNe]�(NNKbKaNNK\K[KZKYKXKWKVKUKTKSKRKQNNNNNNNNNNNNNNNNNNNK/NNNNNNNNK$K#K"K!K KKKNNNNNNNNNNKKKKKKK
K	KKKKKKKKKNNNNNNNNNNNNNNNNNNNe]�(NNKaK`K_K^K]K\K[NNNNNNNNNNNNNNNNNNNNNNNNNNNNK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKNNNNNNNNNNNNNNNNNKKKKKKKKK KNNNNNNNNNNNNNNNNNNNe]�(NNKbKaK`K_K^K]K\NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK#K"K!K KNNNNNNNNNNNNNNNNNK	KKKKKKKKKNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK$K#K"K!K NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK%K$K#K"K!NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeeh:�1A: Sacked Tower�jt9  }�(Kj�  )��}�(j�  KJj�  j�  j�  �Features.Features��Chest���)��}�(hWjײ  h=h>hO]�hj��  h:jڲ  ubjv9  K�ID�Khj��  h:jڲ  ubKj�  )��}�(j�  KGj�  j�  j�  j۲  )��}�(hWj�  h=h>hO]�hj��  h:jڲ  ubjv9  Kj߲  Khj��  h:jڲ  ubKj�  )��}�(j�  KNj�  j�  j�  j  jv9  K	j߲  Khh<h:�Item�ubKj�  )��}�(j�  Kj�  j�  j�  j۲  )��}�(hWj�  h=h>hO]�hj��  h:jڲ  ubjv9  Kj߲  Khj��  h:jڲ  ubKj�  )��}�(j�  Kj�  j�  j�  j۲  )��}�(hWj�  h=h>hO]�hj��  h:jڲ  ubjv9  Kj߲  Khj��  h:jڲ  ubKj�  )��}�(j�  K
j�  j�  j�  jl9  )��}�(hWNh7h5h=]�(K�K�Keh@�h5��coins�Kh�$�h:�
Gold Coins�ubjv9  Kj߲  Khjb  h:�Health�ubK#j�  )��}�(j�  K6j�  j�  j�  jٲ  �Brush���)��}�(hWj��  h=]�(KKnKehj�  h:j��  ubjv9  K#j߲  K#hj�  h:j��  ubK$j�  )��}�(j�  K7j�  j�  j�  j��  )��}�(hWj�  h=j�  hj�  h:j��  ubjv9  K#j߲  K$hj�  h:j��  ubK&j�  )��}�(j�  K8j�  j�  j�  h�jv9  K(j߲  K&hjb  h:j��  ubK'j�  )��}�(j�  KNj�  j�  j�  j۲  )��}�(hWj�  h=h>hO]�hj��  h:jڲ  ubjv9  K(j߲  K'hj��  h:jڲ  ubK*j�  )��}�(j�  KNj�  j�  j�  j۲  )��}�(hWj�  h=h>hO]�hj��  h:jڲ  ubjv9  K)j߲  K*hj��  h:jڲ  ubK,j�  )��}�(j�  K9j�  j�  j�  j۲  )��}�(hWj�  h=h>hO]�hj��  h:jڲ  ubjv9  K+j߲  K,hj��  h:jڲ  ubK.j�  )��}�(j�  Kj�  j�  j�  jn�  )��}�(�
stealthVal�K hK �isAfraid��hKhKh	]�hNh*�h&Kh'K �	cowardice�G?�      �
dropChance�K(j~  Kh(�h)NhKd�
alliesList�]�(j�  j�  )��}�(j�  Kj�  j�  j�  jn�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�      j�  K(j~  Kh(�h)NhKdj �  ]�(j�  j"�  j�  )��}�(j�  Kj�  j�  j�  jn�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�      j�  K(j~  Kh(�h)NhKdj �  ]�(j�  j�  )��}�(j�  Kj�  j�  j�  jn�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�      j�  K(j~  Kh(�h)NhKdj �  ]�(j"�  j.�  j(�  j�  )��}�(j�  Kj�  j�  j�  jn�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�      j�  K(j~  Kh(�h)NhKdj �  ]�(j.�  j(�  j4�  j�  )��}�(j�  Kj�  j�  j�  jd�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�������j�  K(j~  Kh(�h)NhKdj �  ]�(j4�  j�  )��}�(j�  Kj�  j�  j�  jb�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G        j�  K(j~  Kh(�h)NhKdj �  ]�(j@�  j�  )��}�(j�  Kj�  j�  j�  jd�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�������j�  K(j~  Kh(�h)NhKdj �  ]�(j@�  jF�  j:�  eh,�h/j �  )��}�(h5�h&K h6KhXKh7h8h9�hKh:j�  h;�hKhh<h=h>h?�h@�hAK ubhBKhC�hEK hFhc)��}�(h5�h&Kh6Kh7hKh9�hKh:hbh;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNK
hO]�jy  K �hearingDist�KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  ��lastPlayerMap�Nh:�Goblin Lancer�hWjF�  �necklace�N�accuracy�K h=]�(K�KKe�lastPlayerLoc�N�	sightDist�K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  KKj߲  KOhj��  h:�Enemy�ubj:�  eh,�h/j  )��}�(h5�h&K h6KhXKh7hoh9�hKh:j  h;�hKhh<h=h>h?�h@�hAK ubhBKhC�hEK hFh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^j"�  )��}�(h6K7hKh7h^h=h>h?�h@�h5�hXK2hh<h:�Iron Breastplate�ubhj��  j  �jU�  Nh:�Goblin Stonewall�hWj@�  jW�  NjX�  K h=jY�  jZ�  Nj[�  KhXK hVhg)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:hjububjv9  KKj߲  KNhj��  h:j^�  ubjF�  j:�  eh,�h/j �  )��}�(h5�h&K h6KhXKh7h8h9�hKh:j�  h;�hKhh<h=h>h?�h@�hAK ubhBKhC�hEK hFhc)��}�(h5�h&Kh6Kh7hKh9�hKh:hbh;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:jV�  hWj:�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  KNj߲  KRhj��  h:j^�  ubeh,�h/h�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhBKhC�hEK hFh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKub�optionalTargets�]�j�  j�  ��ahL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:�Goblin Thief�hWj4�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  KGj߲  K[hj��  h:j^�  ubeh,�h/h�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhBKhC�hEK hFh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubjy�  ]�j{�  ahL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:j��  hWj.�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  KEj߲  KKhj��  h:j^�  ubj(�  j"�  eh,�h/h�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhBKhC�hEK hFh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubjy�  ]�j{�  ahL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:j��  hWj(�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  KEj߲  KWhj��  h:j^�  ubj4�  eh,�h/h�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhBKhC�hEK hFh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubjy�  ]�j{�  ahL�j{  K hNKhO]�hc)��}�(hWNh5�h&Kh6Kh7hKh9�hKh:hbh;�hKhh<h=h>h?�h@�hKhAKubajy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:j��  hWj"�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  KEj߲  KPhj��  h:j^�  ubeh,�h/h�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhBKhC�hEK hFh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubjy�  ]�j{�  ahL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:j��  hWj�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  KBj߲  K.hj��  h:j^�  ubK/j�  )��}�(j�  Kj�  j�  j�  jb�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G        j�  K(j~  Kh(�h)NhKdj �  ]�j��  ah,�h/j  )��}�(h5�h&K h6KhXKh7hoh9�hKh:j  h;�hKhh<h=h>h?�h@�hAK ubhBKhC�hEK hFh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^j"�  )��}�(h6K7hKh7h^h=h>h?�h@�h5�hXK2hh<h:jg�  ubhj��  j  �jU�  Nh:jh�  hWj��  jW�  NjX�  K h=jY�  jZ�  Nj[�  KhXK hVhg)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:hjububjv9  K,j߲  K/hj��  h:j^�  ubK0j�  )��}�(j�  Kj�  j�  j�  j۲  )��}�(hWj��  h=]�(KQKOKehO]�(jj9  )��}�(�
arrowCount�Kh7h5h=h>h@�h5�h�i�h:�Bundle of Arrows�ubj  )��}�(h5�h&K h6KhXKh7hoh9�hKh:j  h;�hKhh<h=h>h?�h@�hAK ubhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYubjl9  )��}�(h7h5h=j��  h@�h5�j��  Khj��  h:j��  ubehj��  h:jڲ  ubjv9  K,j߲  K0hj��  h:jڲ  ubK1j�  )��}�(j�  K
j�  j�  j�  jf�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G        j�  K(j~  Kh(�h)NhKdj �  ]�(j��  jҳ  j�  )��}�(j�  K
j�  j�  j�  jf�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G        j�  K(j~  Kh(�h)NhKdj �  ]�(j��  jҳ  jس  eh,�h/NhBKhC�hEK hFhH)��}�(h5�h&Kh6Kh7hKh9�hKh:hGh;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:�Goblin Berserker�hWjس  jW�  NjX�  K h=jY�  jZ�  Nj[�  KhXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  K0j߲  K:hj��  h:j^�  ubeh,�h/NhBKhC�hEK hFhH)��}�(h5�h&Kh6Kh7hKh9�hKh:hGh;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNK
hO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:j�  hWjҳ  jW�  NjX�  K h=jY�  jZ�  Nj[�  KhXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  K,j߲  K1hj��  h:j^�  ubK3j�  )��}�(j�  Kj�  j�  j�  jl�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?��Q�j�  K(j~  Kh(�h)NhKdj �  ]�(j�  j�  )��}�(j�  Kj�  j�  j�  jb�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G        j�  K(j~  Kh(�h)NhKdj �  ]�(j�  j��  eh,�h/j  )��}�(h5�h&K h6KhXKh7hoh9�hKh:j  h;�hKhh<h=h>h?�h@�hAK ubhBKhC�hEK hFh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^j"�  )��}�(h6K7hKh7h^h=h>h?�h@�h5�hXK2hh<h:jg�  ubhj��  j  �jU�  Nh:jh�  hWj��  jW�  NjX�  K h=jY�  jZ�  Nj[�  KhXK hVhg)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:hjububjv9  K1j߲  K=hj��  h:j^�  ubj�  )��}�(j�  K!j�  j�  j�  jl�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?��Q�j�  K(j~  Kh(�h)NhKdj �  ]�(j�  j��  j�  eh,�h/NhBKhC�hEK hFhl)��}�(h5�h&Kh6Kh7hoh9�hKh:hkh;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:�Goblin Grunt�hWj�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  K2j߲  K>hj��  h:j^�  ubeh,�h/NhBKhC�hEK hFhl)��}�(h5�h&Kh6Kh7hoh9�hKh:hkh;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:j�  hWj�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  K-j߲  K3hj��  h:j^�  ubK4j�  )��}�(j�  K2j�  j�  j�  hyjv9  K-j߲  K4hh<h:j�  ubK8j�  )��}�(j�  Kj�  j�  j�  h�)��}�(hWj�  h5�h�Kh7h5hK h:h�h�KhKhh�h=h>h�Kh@�h�h�ubjv9  K/j߲  K8hjb  h:j��  ubK9j�  )��}�(j�  Kj�  j�  j�  jn�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�      j�  K(j~  Kh(�h)NhKdj �  ]�(j�  )��}�(j�  Kj�  j�  j�  jl�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?��Q�j�  K(j~  Kh(�h)NhKdj �  ]�(j(�  j�  )��}�(j�  Kj�  j�  j�  jb�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G        j�  K(j~  Kh(�h)NhKdj �  ]�(j(�  j.�  eh,�h/j  )��}�(h5�h&K h6KhXKh7hoh9�hKh:j  h;�hKhh<h=h>h?�h@�hAK ubhBKhC�hEK hFh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^j"�  )��}�(h6K7hKh7h^h=h>h?�h@�h5�hXK2hh<h:jg�  ubhj��  j  �jU�  Nh:jh�  hWj.�  jW�  NjX�  K h=jY�  jZ�  Nj[�  KhXK hVhg)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:hjububjv9  K9j߲  K@hj��  h:j^�  ubj"�  j�  )��}�(j�  Kj�  j�  j�  jn�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�      j�  K(j~  Kh(�h)NhKdj �  ]�(j(�  j.�  j"�  j>�  eh,�h/h�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhBKhC�hEK hFh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubjy�  ]�j{�  ahL�j{  K hNK	hO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:j��  hWj>�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  K>j߲  KBhj��  h:j^�  ubeh,�h/NhBKhC�hEK hFhl)��}�(h5�h&Kh6Kh7hoh9�hKh:hkh;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:j�  hWj(�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  K9j߲  K?hj��  h:j^�  ubj.�  j"�  j>�  eh,�h/h�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhBKhC�hEK hFh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubjy�  ]�j{�  ahL�j{  K hNKhO]�h[)��}�(h6KhKh7h^hWNh=h>h?�h@�h5�hXKhh<h:h_ubajy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:j��  hWj"�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  K?j߲  K9hj��  h:j^�  ubK:jس  K<j�  )��}�(j�  Kj�  j�  j�  j]�  jv9  K1j߲  K<hh<h:j�  ubK=j��  K>j�  K?j(�  K@j.�  KBj>�  KCj�  )��}�(j�  Kj�  j�  j�  jh�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�      j�  K(j~  Kh(�h)NhKdj �  ]�(jf�  j�  )��}�(j�  Kj�  j�  j�  jl�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?��Q�j�  K(j~  Kh(�h)NhKdj �  ]�(jf�  jl�  j�  )��}�(j�  Kj�  j�  j�  jh�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�      j�  K(j~  Kh(�h)NhKdj �  ]�(jf�  jl�  jr�  eh,�h/NhBKhC�hEKhFh�)��}�(h5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:�Goblin Archer�hWjr�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K
hXK hVhx)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:h{ububjv9  K?j߲  KLhj��  h:j^�  ubeh,�h/NhBKhC�hEK hFhl)��}�(h5�h&Kh6Kh7hoh9�hKh:hkh;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:j�  hWjl�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  K=j߲  KHhj��  h:j^�  ubjr�  eh,�h/NhBKhC�hEKhFh�)��}�(h5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:j~�  hWjf�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K
hXK hVhx)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:h{ububjv9  K:j߲  KChj��  h:j^�  ubKDj�  )��}�(j�  KLj�  j�  j�  j۲  )��}�(hWj��  h=h>hO]�hj��  h:jڲ  ubjv9  K;j߲  KDhj��  h:jڲ  ubKEj�  )��}�(j�  K9j�  j�  j�  �Features.Stairs��StairUp���)��}�(j�  K9j�  j�  hWj��  j�  Njv9  K<j߲  J�����moveCost�Kh:�Stairs�ubjv9  K<j߲  KEhj5�  h:�	Stairs Up�ubKFj�  KGj�  )��}�(j�  K5j�  j�  j�  jn�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�      j�  K(j~  Kh(�h)NhKdj �  ]�j��  ah,�h/h�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhBKhC�hEK hFh�)��}�(h5�h&Kh6Kh7hoh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubjy�  ]�j{�  ahL�j{  K hNK
hO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK\K[KZKYNNNNNNNNNNNNNNNNNKGKHKIKJKKKLNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK[KZKYKXNNNNNNNNNNNNNNNNNKFKGKHKIKJKKNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�KNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK\K[KZKYKXKWNNNNNNNNNNNNNNNNNKEKFKGKHKIKJNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�KK~K}K|K{KzKyKxKwKvKuNNNNNNNNNNNNNNNNNNNKaK`K_K^K]K\K[KZKYKXKWKVNNNNNNNNNNNNNNNNNKDKEKFKGKHKIKJKKKLNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�KNNNNNNNNKtNNNNNNNNNNNNNNNNNNNKbNNNNNKZKYKXKWKVKUNNNNNNNNNNNNNNNNNKCKDKEKFKGKHKIKJKKNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNKsNNNNNNNNNNNNNNNNNNNKcNNNNNKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJNNNNNNNKBKCKDKEKFKGKHKIKJNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNKrNNNNKmKlKkKjKkKlNNNNNNNNNKdNNNNNKZNNNNNNNNNNNNNNKIKHKGKFKEKDKCKBKAKBKCKDKEKFKGKHKINNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNKqKpKoKnKmKlKkKjKiKjKkKlKmKlKkKjKiKhKgKfKeNNNNNK[NNNNNNNNNNNNNNNNNNNNNNK@KAKBKCKDKEKFKGKHNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNKkKjKiKhNNNNNNNNNNNNNNNNNKZNNNNNNNNNNNNNNNNNNNNNNK?NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNKjKiKhKgNNNNNNNNNNNNNNNNNKYNNNNNNNNNNNNNNNNNNNNNNK>NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNKiKhKgKfKgKhNNNNNNNNNNNNNNNKXNNNNNNNNNNNNNNNNNNNNNNK=NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNKhKgKfKeKfKgNNNNNNNNNNNNNNNKWNNNNNNNNNNNNNNNNNNNNNNK<NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNKgKfKeKdKeKfNNNNNNNNNNNNNNNKVNNNNNNNNNNNNNNNNNNNNNNK;NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNKfKeKdKcKdKeNNNNNNNNNNNNNNNKUNNNNNNNNNNNNNNNNNNNNNNK:NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNKbNNNNNNNNNNNNNNNNNKTKSKRKQKPKOKNNNNNNNNNNNNNNNNNK9NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNKaNNNNNNNNNNNNNNNNNNNNNNNKMNNNNNNNNNNNNNNNNK8NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNK`NNNNNNNNNNNNNNNNNNNNNNNKLNNNNNNNNNNNNNNNNK7NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNK_K^NNNNNNNNNNNNNNNNNNNNNNKKNNNNNNNNNNNNNNNNK6K5K4NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNK]NNNNNNNNNNNNNNNNNNNNNNKJNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�K�K�K�NNNNNNNNNNNNNNNNNNNNNK\NNNNNNNNNNNNNNNNNNNNNNKINNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNKaK`K_K^K]K\K[KZKYKXNNNNNNNNNNNNNNNNNNNKHNNNNNNNNNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKONNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNK0NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNKaK`K_K^K]K\K[KZKYKXNNNNNNNKNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNK/NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNKbKaK`NNNNK[KZKYNNNNNNNKMNNNNNNNNNNNKENNNNNNNNNNNNNNNNK0K/K.K-K,K-K.K/K0K1NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNKcKbKaNNNNK\K[KZNNNNNNNKLNNNNNNNNKCKBKCKDKEKFKGKHKGNNNNNNNNK2K1K0K/K.K-K,K+K,K-K.K/K0NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�KNNNNNNNNKjKiKhKgKfKeKdKcKbNNNNK]K\K[NNNNNNNKKNNNNNNNNKBKAKBKCKDKEKFKGKFNNNNNNNNK3NNK.K-K,K+K*K+K,K-K.K/NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�KK~NNNNNNNNKkNNNNNKeKdKcNNNNK^K]K\NNNNNNNKJKIKHKGKFKEKDKCKBKAK@KAKBKCKDKEKFKENNNNNNNNK4NNK-K,K+K*K)K*K+K,K-K.NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�KK~K}NNNNNNNNKlNNNNNKfKeKdKcKbKaK`K_K^K]NNNNNNNNNNNNNNNNK@K?K@KAKBKCKDKEKDNNNNNNNNK5NNNNK*K)K(K)K*K+K,K-NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK}K|NNNNNNNNKmNNNNNKgKfKeKdKcKbKaK`K_K^NNNNNNNNNNNNNNNNK?K>K?K@KAKBKCKDKCNNNNNNNNK6NNNNK)K(K'K(K)K*K+K,NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK|K{NNNNNNNNKnNNNNNNKgNNNNNNNNNNNNNNNNNNNNNNNNK>K=K>K?K@KAKBKCKBNNNNNNNNK7NNNNNNK&NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK{KzNNNNNNNNKoNNNNNNKhNNNNNNNNNNNNNNNNNNNNNNNNK=K<K=K>K?K@KAKBKAK@K?K>K=K<K;K:K9K8NNNNNNK%NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNKzKyKxKwKvKuKtKsKrKqKpNNNNNNKiNNNNNNNNNNNNNNNNNNNNNNNNNK;NNNNNNNNNNNNNNNNNNNNNNK$K#K"K!K NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK{NNNNNNNNNNNNNNNNKjNNNNNNNNNNNNNNNNNNNNNNNNNK:NNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK|NNNNNNNNNNNNNNNNKkNNNNNNNNNNNNNNNNNNNNNNNNNK9K8K7K6K5NNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK}NNNNNNNNNNNNNNNNKlNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�K�K�K�KK~NNNNNNNNNNNNNNNNKmNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNNKnNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNNKoNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNNKpNNNNNNNNNNNNNNNNNNNNNNNK2K1K0K/K.K/K0K1K0NNNNNNNNNNNNNNNNNNKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNNKqNNNNNNNNNNNNNNNNNNNNNNNK1K0K/K.K-K.K/K0K/NNNNNNNNNNNNNNNNNNKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNKsKrKsKtKuKvKwKxKyNNNNNNNNNNNNNNNNK0K/K.K-K,K-K.K/K.NNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNKzKyKxKwKvKuKtKsKtKuKvKwKxKyKzNNNNNNNNNNNNNNNNK/K.K-K,K+K,K-K.K-NNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK{NNNNNKuKtKuKvKwKxKyKzK{NNNNNNNNNNNNNNNNK.K-K,K+K*K+K,K-K,NNNNNNNNNK KKKKKKKKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK|NNNNNKvKuKvKwKxKyKzK{K|NNNNNNNNNNNNNNNNK-K,K+K*K)K*K+K,K+K*K)K(K'K&K%K$K#K"K!NNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK}NNNNNKwKvKwKvKwKxKyKzK{NNNNNNNNNNNNNNNNK,K+K*K)K(K)K*K+K,NNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNK�K�K�K�NNNNNNNNK~NNNNNKxKwKvKuKvKwKxKyKzNNNNNNNNNNNNNNNNK+K*K)K(K'K(K)K*K+NNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNK�K�K�K�NNNNNNNNKNNNNNKwKvKuKtKuKvKwKxKyNNNNNNNNNNNNNNNNK*K)K(K'K&K'K(K)K*NNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK�NNNNNKvKuKtKsKtKuKvKwKxNNNNNNNNNNNNNNNNK)K(K'K&K%K&K'K(K)NNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK�NNNNNKuKtKsKrKsKtKuKvKwNNNNNNNNNNNNNNNNNNNNK$NNNNNNNNNNNNNNNKKKKKK	K
KKKKNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�NNNNNKtKsKrKqKrKsKtKuKvNNNNNNNNNNNNNNNNNNNNK#NNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNNNNKpNNNNNNNNNNNNNNNNNNNNNNNNNK"NNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�K�K�K�K�NNNNNNNNNNNNNNNNNNNKoNNNNNNNNNNNNNNNNNNNNNNNNNK!K KKKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNK�NNNNNNNNNNNNNNNNNNNKnNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNK NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKNNNNNNNNNNNNNNNNNNNKmKlKkKjKiNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�KK~K}K|K{NNNNNNNNNNNNNNNNNNNNKhNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�KK~K}K|K{KzNNNNNNNNNNNNNNNNNNNNKgNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNKKKKKKKK	K
NNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�KK~K}K|K{KzKyKxKwKvKuKtKsKrKqNNNNNNNNNKgKfKeKfKgNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNKKKKKKK	K
KNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�KK~K}K|K{KzNNNNNNNKpNNNNNNNNNKfKeKdKeKfNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNKKKKKK	K
KKNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�KNNNK{NNNNNNNKoNNNNNNNKgKfKeKdKcKdKeNNNNNNNNNNNNNNNNNNKKKKKKKKKKKKKKKNNKKKKK	K
KKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�NNNK|NNNNNNNKnNNNNNNNKfKeKdKcKbKcKdNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNKNNKKKK	K
KKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�NNNK}NNNNNNNKmKlKkKjKiKhKgKfKeKdKcKbKaKbKcNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNKKK
K	KK	K
KKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�KK~NNNNNNNNNNNNNNNKdKcKbKaK`KaKbNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNK
K	K
KKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNNNKcKbKaK`K_K`KaNNNNNNNNNNNNNNNNNNK KKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNK^NNNNNNNNNNNNNNNNNNNNK!K KKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNK]NNNNNNNNNNNNNNNNNNNNK"K!K KKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNK\NNNNNNNNNNNNNNNNNNNNK#K"K!K KKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNK[NNNNNNNNNNNNNNNNNNNNK$K#K"K!K KKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNK�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNNKZNNNNNNNNNNNNNNNNNNNNNK$NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNKYNNNNNNNNNNNNNNNNNNNNNK%NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNK~NNNNNNNNNNNNNNNNNNNNNNNNNKVKWKXNNNNNNNNNNNNNNNNNNNNNK&NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNK}NNNNNNNNNNNNNNNNNNNNNNNNNKUNNNNNNNNNNNNNNNNNNNNNNNK'NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNK|NNNNNNNNNNNNNNNNNNNNNNNNNKTNNNNNNNNNNNNNNNNNK.K-K,K+K*K)K(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNK{NNNNNNNNNNNNNNNNNNNNNKWKVKUKTKSKRKQKPNNNNNNNNNNNNNNK/NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK{KzKyKxKwKvKuNNNNNNNNNNNNNNNNKVKUKTKSKRKQKPKOKNKMKLKKKJNNNNNNNNNK0NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKzKyKxKwKvKuKtNNNNNNNNNNNNNNNNKWKVKUKTKSKRKQKPNNNNKINNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKyKxKwKvKuKtKsNNNNNNNNNNNNNNNNKXKWNNNKSKRKQNNNNKHNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKxKwKvKuKtKsKrNNNNNNNNNNNNNNNNKYKXNNNKTKSKRNNNNKGNNNNNNNNK4K3K4K5K6K7K8K9NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKwKvKuKtKsKrKqNNNNNNNNNNNNNNNNKZKYNNNKUKTKSNNNNKFNNNNNNNNK5K4K5K6K7K8K9K:NNNNNNNNNNNNNNNNNKRKSKTKUKVKWKXKYKZK[NNNNNNNNNNNNNNNNNNNe]�(NNKvKuKtKsKrKqKpNNNNNNNNKcKbKaK`K_K^K]K\K[KZKYKXKWKVKUKTNNNNKENNNNNNNNK6K5K6K7K8K9K:K;NNNNNNNNNNNNNNNNNKQKRKSKTKUKVKWKXKYKZNNNNNNNNNNNNNNNNNNNe]�(NNKwKvNNKqKpKoNNNNNNNNKdNNNNNNNK\K[KZKYKXKWKVKUNNNNKDNNNNNNNNK7K6K7K8K9K:K;K<K=K>K?K@KAKBKCKDKEKFKGNNNNNNKPKQKRKSKTKUKVKWKXKYNNNNNNNNNNNNNNNNNNNe]�(NNKvKuNNKpKoKnKmKlKkKjKiKhKgKfKeNNNNNNNNNNNNNNNNNNNKCNNNNNNNNK8K7K8K9K:K;K<K=NNNNNNNNNNKHKIKJKKKLKMKNKOKPKQKRKSKTKUKVKWKXNNNNNNNNNNNNNNNNNNNe]�(NNKuKtKsKrKqKpKoNNNNNNNNNNNNNNNNNNNNNNNNNNNNKBKAK@K?K>K=K<K;K:K9K8K9K:K;K<K=K>NNNNNNNNNNNNNNNNNKPKQKRKSKTKUKVKWKXKYNNNNNNNNNNNNNNNNNNNe]�(NNKvKuKtKsKrKqKpNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK;K<K=K>K?NNNNNNNNNNNNNNNNNKQKRKSKTKUKVKWKXKYKZNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK<K=K>K?K@NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK=K>K?K@KANNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeeh:j��  hWj��  jW�  NjX�  K h=jY�  jZ�  ]�(K6KFej[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  Kj߲  KGhj��  h:j^�  ubKHjl�  KKj.�  KLjr�  KMj�  )��}�(j�  Kj�  j�  j�  jh�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�      j�  K(j~  Kh(�h)NhKdj �  ]�j�  ah,�h/NhBKhC�hEKhFh�)��}�(h5�h&Kh6Kh7hKh9�hKh:h�h;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:j~�  hWj�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K
hXK hVhx)��}�(h6KhKh7hVh=h>h?�h@�h5�hXKhh<h:h{ububjv9  KJj߲  KMhj��  h:j^�  ubKNj@�  KOjF�  KPj"�  KQj�  )��}�(j�  Kj�  j�  j�  j۲  )��}�(hWj%�  h=jų  hO]�(jl9  )��}�(h7h5h=j��  h@�h5�j��  Khj��  h:j��  ubh�)��}�(hKh7h�h=h>h@�h5�hh�h�hh:h�ubj�  )��}�(h5�h&Kh6Kh7hKh9�hKh:j�  h;�hKhh<h=h>h?�h@�hKhAKubjl9  )��}�(h7h5h=j��  h@�h5�j��  Khj��  h:j��  ubehj��  h:jڲ  ubjv9  KMj߲  KQhj��  h:jڲ  ubKRj:�  KSj�  )��}�(j�  Kj�  j�  j�  j۲  )��}�(hWj2�  h=jų  hO]�(h�)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h�ubhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYubj_  )��}�(h7h5h=h>h@�h5�hjb  jc  Kh:jd  ubjl9  )��}�(h7h5h=j��  h@�h5�j��  Khj��  h:j��  ubehj��  h:jڲ  ubjv9  KNj߲  KShj��  h:jڲ  ubKTj�  )��}�(j�  Kj�  j�  j�  jd�  )��}�(j�  K hK j�  �hKhKh	]�hNh*�h&Kh'K j�  G?�������j�  K(j~  Kh(�h)NhKdj �  ]�j?�  ah,�h/j �  )��}�(h5�h&K h6KhXKh7h8h9�hKh:j�  h;�hKhh<h=h>h?�h@�hAK ubhBKhC�hEK hFhc)��}�(h5�h&Kh6Kh7hKh9�hKh:hbh;�hKhh<h=h>h?�h@�hKhAKubhL�j{  K hNKhO]�jy  K jQ�  KhMKj|  ]�h^h[)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h_ubhj��  j  �jU�  Nh:jV�  hWj?�  jW�  NjX�  K h=jY�  jZ�  Nj[�  K	hXK hVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYububjv9  KOj߲  KThj��  h:j^�  ubKVj�  )��}�(j�  KLj�  j�  j�  j۲  )��}�(hWjO�  h=jų  hO]�(hS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYubj�  )��}�(h5�h&Kh6Kh7hKh9�hKh:j�  h;�hKhh<h=h>h?�h@�hKhAKubh�)��}�(h5�h��50      Kh7h5hK h:h�h�KhKhh�h=h>h�Kh@�h�h�ubjl9  )��}�(h7h5h=j��  h@�h5�j��  Khj��  h:j��  ubehj��  h:jڲ  ubjv9  KOj߲  KVhj��  h:jڲ  ubKWj(�  KXj�  )��}�(j�  Kj�  j�  j�  j��  )��}�(hWj\�  h=j�  hj�  h:j��  ubjv9  KPj߲  KXhj�  h:j��  ubKYj�  )��}�(j�  Kj�  j�  j�  j��  )��}�(hWj`�  h=j�  hj�  h:j��  ubjv9  KPj߲  KYhj�  h:j��  ubKZj�  )��}�(j�  Kj�  j�  j�  j��  )��}�(hWjd�  h=j�  hj�  h:j��  ubjv9  KPj߲  KZhj�  h:j��  ubK[j4�  K]j�  )��}�(j�  Kj�  j�  j�  j��  )��}�(hWjh�  h=j�  hj�  h:j��  ubjv9  KQj߲  K]hj�  h:j��  ubKbj�  )��}�(j�  Kj�  j�  j�  j��  )��}�(hWjl�  h=j�  hj�  h:j��  ubjv9  KRj߲  Kbhj�  h:j��  ubKcj�  )��}�(j�  Kj�  j�  j�  j��  )��}�(hWjp�  h=j�  hj�  h:j��  ubjv9  KRj߲  Kchj�  h:j��  ubKdj�  )��}�(j�  Kj�  j�  j�  j��  )��}�(hWjt�  h=j�  hj�  h:j��  ubjv9  KRj߲  Kdhj�  h:j��  ubKfj�  )��}�(j�  KPj�  j�  j�  j �  )��}�(hWj�  )��}�(j�  KFj�  j�  j�  jz�  jv9  KRj߲  K�hh<h:j�  ubh5�h&K h6KhXKh7h8h9�hKh:j�  h;�hKhh<h=h>h?�h@�hAK ubjv9  KRj߲  Kfhh<h:j�  ubKhj�  )��}�(j�  KOj�  j�  j�  j��  �	StairDown���)��}�(j�  KOj�  j�  hWj~�  j�  Njv9  KSj߲  J����h:j��  j��  Kubjv9  KSj߲  KhhjM�  h:�Stairs Down�ubKij�  )��}�(j�  Kj�  j�  j�  j��  jv9  KTj߲  Kihh<h:j�  ubKjj�  )��}�(j�  K6j�  j�  j�  hTjv9  K3j߲  Kjhh<h:hYubKkj�  )��}�(j�  K6j�  j�  j�  hdjv9  K3j߲  Kkhh<h:hbubKlj�  )��}�(j�  K6j�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  K3j߲  Klhj��  h:j��  ubKmj�  )��}�(j�  K6j�  j�  j�  hTjv9  K3j߲  Kmhh<h:hYubKnj�  )��}�(j�  K6j�  j�  j�  h\jv9  K3j߲  Knhh<h:h_ubKoj�  )��}�(j�  K6j�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  K3j߲  Kohj��  h:j��  ubKpj�  )��}�(j�  K6j�  j�  j�  hdjv9  K3j߲  Kphh<h:hbubKqj�  )��}�(j�  K6j�  j�  j�  h`jv9  K3j߲  Kqhh<h:h_ubKrj�  )��}�(j�  K6j�  j�  j�  jj9  )��}�(jɳ  Kh7h5hWNh=h>h@�h5�hjʳ  h:j˳  ubjv9  K3j߲  Krhjʳ  h:j˳  ubKsj�  )��}�(j�  K6j�  j�  j�  hdjv9  K3j߲  Kshh<h:hbubKtj�  )��}�(j�  K6j�  j�  j�  hpjv9  K3j߲  Kthh<h:h_ubKuj�  )��}�(j�  K6j�  j�  j�  htjv9  K3j߲  Kuhh<h:hvubKvj�  )��}�(j�  K6j�  j�  j�  hhjv9  K2j߲  Kvhh<h:hjubKwj�  )��}�(j�  K6j�  j�  j�  hmjv9  K2j߲  Kwhh<h:hkubKxj�  )��}�(j�  K6j�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  K2j߲  Kxhj��  h:j��  ubKyj�  )��}�(j�  K4j�  j�  j�  h�jv9  K!j߲  Kyhh<h:hjubKzj�  )��}�(j�  K4j�  j�  j�  h�jv9  K!j߲  Kzhh<h:hkubK{j�  )��}�(j�  K4j�  j�  j�  jj9  )��}�(jɳ  Kh7h5hWNh=h>h@�h5�hjʳ  h:j˳  ubjv9  K!j߲  K{hjʳ  h:j˳  ubK|j�  )��}�(j�  K4j�  j�  j�  h�jv9  Kj߲  K|hh<h:h{ubK}j�  )��}�(j�  K4j�  j�  j�  h�jv9  Kj߲  K}hh<h:h�ubK~j�  )��}�(j�  K4j�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K~hj��  h:j��  ubKj�  )��}�(j�  K5j�  j�  j�  h�jv9  Kj߲  Khh<h:h{ubK�j�  )��}�(j�  K5j�  j�  j�  h�jv9  Kj߲  K�hh<h:h�ubK�j�  )��}�(j�  K5j�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  K!j�  j�  j�  h�jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  K!j�  j�  j�  h�jv9  Kj߲  K�hh<h:hkubK�j�  )��}�(j�  K!j�  j�  j�  h�jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  K!j�  j�  j�  h�jv9  Kj߲  K�hh<h:h_ubK�j�  )��}�(j�  K!j�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  K j�  j�  j�  h�jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  K j�  j�  j�  h�jv9  Kj߲  K�hh<h:hGubK�j�  )��}�(j�  K j�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:hbubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh�h:h�ubK�j�  )��}�(j�  K
j�  j�  j�  h�jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  K
j�  j�  j�  h�jv9  Kj߲  K�hh<h:hGubK�j�  )��}�(j�  K
j�  j�  j�  h�jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  K
j�  j�  j�  h�jv9  Kj߲  K�hh<h:h_ubK�j�  )��}�(j�  K
j�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:hbubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:h_ubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:hvubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:h{ubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:h�ubK�j�  )��}�(j�  K	j�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:hbubK�j�  )��}�(j�  K	j�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:hjubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:h�ubK�j�  )��}�(j�  K	j�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:h{ubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:h�ubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:hjubK�j�  )��}�(j�  K	j�  j�  j�  h�jv9  Kj߲  K�hh<h:h�ubK�j�  )��}�(j�  K	j�  j�  j�  jj9  )��}�(jɳ  Kh7h5hWNh=h>h@�h5�hjʳ  h:j˳  ubjv9  Kj߲  K�hjʳ  h:j˳  ubK�j�  )��}�(j�  Kj�  j�  j�  h�jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  Kj�  j�  j�  h�jv9  Kj߲  K�hh<h:h�ubK�j�  )��}�(j�  Kj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  Kj�  j�  j�  h�jv9  K	j߲  K�hh<h:hYubK�j�  )��}�(j�  Kj�  j�  j�  h�jv9  K	j߲  K�hh<h:hGubK�j�  )��}�(j�  Kj�  j�  j�  h�jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  Kj�  j�  j�  h�jv9  Kj߲  K�hh<h:hbubK�j�  )��}�(j�  Kj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  K/j�  j�  j�  h�jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  K/j�  j�  j�  h�jv9  Kj߲  K�hh<h:hkubK�j�  )��}�(j�  K3j�  j�  j�  h�jv9  Kj߲  K�hh<h:h{ubK�j�  )��}�(j�  K3j�  j�  j�  h�jv9  Kj߲  K�hh<h:h�ubK�j�  )��}�(j�  K3j�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  KGj�  j�  j�  h�jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  KGj�  j�  j�  h�jv9  Kj߲  K�hh<h:hkubK�j�  )��}�(j�  KHj�  j�  j�  j  jv9  Kj߲  K�hh<h:h{ubK�j�  )��}�(j�  KHj�  j�  j�  j  jv9  Kj߲  K�hh<h:h�ubK�j�  )��}�(j�  KKj�  j�  j�  j  jv9  Kj߲  K�hh<h:h{ubK�j�  )��}�(j�  KKj�  j�  j�  j  jv9  Kj߲  K�hh<h:h�ubK�j�  )��}�(j�  KKj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  KOj�  j�  j�  j  jv9  Kj߲  K�hh<h:h{ubK�j�  )��}�(j�  KOj�  j�  j�  j  jv9  Kj߲  K�hh<h:h�ubK�j�  )��}�(j�  KOj�  j�  j�  jj9  )��}�(jɳ  Kh7h5hWNh=h>h@�h5�hjʳ  h:j˳  ubjv9  Kj߲  K�hjʳ  h:j˳  ubK�j�  )��}�(j�  KOj�  j�  j�  j  jv9  K	j߲  K�hh<h:j  ubK�j�  )��}�(j�  KOj�  j�  j�  j  jv9  K	j߲  K�hh<h:h_ubK�j�  )��}�(j�  KOj�  j�  j�  j  jv9  K	j߲  K�hh<h:h�ubK�j�  )��}�(j�  KGj�  j�  j�  j  jv9  K
j߲  K�hh<h:hYubK�j�  )��}�(j�  KGj�  j�  j�  j&  jv9  K
j߲  K�hh<h:hGubK�j�  )��}�(j�  KGj�  j�  j�  j  jv9  Kj߲  K�hh<h:hjubK�j�  )��}�(j�  KGj�  j�  j�  j$  jv9  Kj߲  K�hh<h:h�ubK�j�  )��}�(j�  KGj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  KGj�  j�  j�  j   jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  KGj�  j�  j�  j"  jv9  Kj߲  K�hh<h:hkubK�j�  )��}�(j�  KGj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  KHj�  j�  j�  j(  jv9  Kj߲  K�hh<h:hYubK�j�  )��}�(j�  KHj�  j�  j�  j*  jv9  Kj߲  K�hh<h:h�ubK�j�  )��}�(j�  KHj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  Kj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  KNj�  j�  j�  j>  jv9  K'j߲  K�hh<h:h{ubK�j�  )��}�(j�  KNj�  j�  j�  j@  jv9  K'j߲  K�hh<h:h�ubK�j�  )��}�(j�  KNj�  j�  j�  jl9  )��}�(hWjs�  h7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  K'j߲  K�hj��  h:j��  ubK�j�  )��}�(j�  KOj�  j�  j�  j,  jv9  K(j߲  K�hh<h:hYubK�j�  )��}�(j�  KOj�  j�  j�  j0  jv9  K(j߲  K�hh<h:hbubK�j�  )��}�(j�  KOj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  K
hj��  h:j��  ubjv9  K(j߲  K�hj��  h:j��  ubK�j�  )��}�(j�  KOj�  j�  j�  j.  jv9  K)j߲  K�hh<h:hYubK�j�  )��}�(j�  KOj�  j�  j�  j2  jv9  K)j߲  K�hh<h:hbubK�j�  )��}�(j�  KOj�  j�  j�  j<  jv9  K)j߲  K�hh�h:h�ubK�j�  )��}�(j�  KOj�  j�  j�  j4  jv9  K*j߲  K�hh<h:hYubK�j�  )��}�(j�  KOj�  j�  j�  j8  jv9  K*j߲  K�hh<h:hbubK�j�  )��}�(j�  KOj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  K*j߲  K�hj��  h:j��  ubK�j�  )��}�(j�  KNj�  j�  j�  j6  jv9  K*j߲  K�hh<h:h{ubK�j�  )��}�(j�  KNj�  j�  j�  j:  jv9  K*j߲  K�hh<h:h�ubK�j�  )��}�(j�  KNj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  K*j߲  K�hj��  h:j��  ubK�j�  )��}�(j�  KFj�  j�  j�  jT  jv9  K6j߲  K�hh<h:hjubK�j�  )��}�(j�  KFj�  j�  j�  jN  jv9  K6j߲  K�hh<h:h�ubK�j�  )��}�(j�  KFj�  j�  j�  jP  jv9  K6j߲  K�hh�h:h�ubK�j�  )��}�(j�  KFj�  j�  j�  jT  jv9  K6j߲  K�hh<h:hjubK�j�  )��}�(j�  KFj�  j�  j�  jR  jv9  K6j߲  K�hh<h:h_ubK�j�  )��}�(j�  KFj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  K6j߲  K�hj��  h:j��  ubK�j�  )��}�(j�  KFj�  j�  j�  jT  jv9  K6j߲  K�hh<h:hjubK�j�  )��}�(j�  KFj�  j�  j�  jV  jv9  K6j߲  K�hh<h:h_ubK�j�  )��}�(j�  KFj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  K	hj��  h:j��  ubjv9  K6j߲  K�hj��  h:j��  ubK�j�  )��}�(j�  K/j�  j�  j�  je  jv9  KKj߲  K�hh<h:hYubK�j�  )��}�(j�  K/j�  j�  j�  j\  jv9  KKj߲  K�hh<h:hbubK�j�  )��}�(j�  K/j�  j�  j�  j`  jv9  KKj߲  K�hjb  h:jd  ubK�j�  )��}�(j�  K/j�  j�  j�  je  jv9  KKj߲  K�hh<h:hYubK�j�  )��}�(j�  K/j�  j�  j�  jm  jv9  KKj߲  K�hh<h:h_ubK�j�  )��}�(j�  K/j�  j�  j�  jq  jv9  KKj߲  K�hh�h:h�ubK�j�  )��}�(j�  K/j�  j�  j�  jg  jv9  KLj߲  K�hh<h:hYubK�j�  )��}�(j�  K/j�  j�  j�  jk  jv9  KLj߲  K�hh<h:hGubK�j�  )��}�(j�  K/j�  j�  j�  ji  jv9  KMj߲  K�hh<h:hYubK�j�  )��}�(j�  K/j�  j�  j�  jo  jv9  KMj߲  K�hh<h:hGubK�j�  )��}�(j�  KCj�  j�  j�  ju  jv9  KRj߲  K�hh<h:hjubK�j�  )��}�(j�  KCj�  j�  j�  js  jv9  KRj߲  K�hh<h:h�ubK�j�  )��}�(j�  KCj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  KRj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  KCj�  j�  j�  ju  jv9  KRj߲  K�hh<h:hjubK�j�  )��}�(j�  KCj�  j�  j�  h[)��}�(h6KhKh7h^hWjɶ  h=h>h?�h@�h5�hXKhh<h:h_ubjv9  KRj߲  K�hh<h:h_ubK�j�  )��}�(j�  KCj�  j�  j�  jl9  )��}�(hWjͶ  h7h5h=j��  h@�h5�j��  K
hj��  h:j��  ubjv9  KRj߲  K�hj��  h:j��  ubK�j�  )��}�(j�  KFj�  j�  j�  hx)��}�(h6KhKh7hVhWNh=h>h?�h@�h5�hXKhh<h:h{ubjv9  KRj߲  K�hh<h:h{ubK�j�  )��}�(j�  KFj�  j�  j�  jw  jv9  KRj߲  K�hh<h:h�ubK�j�  )��}�(j�  KFj�  j�  j�  jl9  )��}�(hWNh7h5h=j��  h@�h5�j��  Khj��  h:j��  ubjv9  KRj߲  K�hj��  h:j��  ubK�j|�  K�j�  )��}�(j�  KFj�  j�  j�  hS)��}�(h6KhKh7hVhWj۶  h=h>h?�h@�h5�hXK
hh<h:hYubjv9  KRj߲  K�hh<h:hYubK�j�  )��}�(j�  KFj�  j�  j�  hl)��}�(hWj߶  h5�h&Kh6Kh7hoh9�hKh:hkh;�hKhh<h=h>h?�h@�hKhAKubjv9  KRj߲  K�hh<h:hkubu�args�]�(KKe�	equipList�]�(j�  j  j �  hshlhHh�hch�h�hxh[hSj"�  hghh�e�	tilesSeen�]��inSeed�J�x �cLevel�Kubj�  hjv9  KRj߲  KFh:h ubjW�  NjX�  K h=]�(KKYK�e�rightScroll�N�healthCurve�G?�333333j[�  K�Class��Player_Classes��
Spellsword���h^h�)��}�(h6KhKh7h^h=h>h?�h@�h5�hXKhh<h:h�ubhVhS)��}�(h6KhKh7hVh=h>h?�h@�h5�hXK
hh<h:hYubub.