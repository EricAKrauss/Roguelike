��      �__main__��Game���)��}�(�loadRequest���	thePlayer��Player�h��)��}�(�char��@��armorPen�K �range�K�level�K�
hitEffects�]��leftRing�N�recalcTimer�K �expNext�K��skills�}�(�3��	Abilities��Fireball����2�h�Shocking_Grasp����7�h�Ready_for_Battle����4�h�Lightning_Bolt����6�h�Rending_Blow����5�h�Block����1�h�Charge���u�power�K�dodge�K �visible���	rightRing�N�canMove���	recalcMax�K �
countering���
prevTarget�N�skillPoints�K�leftHand��Items.Weapons��Tome���)��}�(�
consumable��h-K �weight�K�type��0H��addPower��hK�name�h8�
usesArrows��hKh�?��color�]�(K�K�K�e�	throwable���
equippable��hK �magPower�Kub�health�K1�blocking���
leftScroll�N�arrows�K�	rightHand�h7�
Greatsword���)��}�(h<�h-Kh=Kh>�2H�h@�hKhAhNhB�hKhhChDhEhF�hG�hKhHKub�invertColor���
initiative�K�gold�MS�items�]�(�Items.Armors��Leather_Helm���)��}�(h=KhKh>�helmet��pObject�NhDhEhF�hG�h<��armorVal�K
hhChA�Leather Helm�ubhX�Leather_Shirt���)��}�(h=KhKh>�armor�h^NhDhEhF�hG�h<�h_KhhChA�Leather Shirt�ubhb)��}�(h=KhKh>heh^NhDhEhF�hG�h<�h_KhhChAhfubh7�Spear���)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhihB�hKhhChDhEhF�hG�hKhHKubhX�	Iron_Helm���)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChA�	Iron Helm�ubh7�	Longsword���)��}�(h^Nh<�h-Kh=Kh>�1H�h@�hKhAhrhB�hKhhChDhEhF�hG�hKhHKubhb)��}�(h=KhKh>heh^NhDhEhF�hG�h<�h_KhhChAhfubh7�Wooden_Shield���)��}�(h^Nh<�h-K h=Kh_Kh>hvh@�hKhA�Wooden Shield�hB�hKhhChDhEhF�hG�hHK ubhX�	Cloth_Hat���)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChA�	Cloth Hat�ubh)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAh�ubhX�Chain_Shirt���)��}�(h=K#hKh>hehDhEhF�hG�h<�h_K#hhChA�Chain Shirt�ub�Items.Consumables��Scroll_of_Fireball���)��}�(h^NhKh>�scroll�hDhEhG�h<�h�s��spell�hhA�Scroll of Fireball�ubhn)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAhqubh)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAh�ubh)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAh�ubh7�Bow���)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubh�)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhs)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAhrhB�hKhhChDhEhF�hG�hKhHKubhs)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAhrhB�hKhhChDhEhF�hG�hKhHKubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhb)��}�(h=KhKh>heh^NhDhEhF�hG�h<�h_KhhChAhfubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhO)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhNhB�hKhhChDhEhF�hG�hKhHKubhn)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAhqubhb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhO)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhNhB�hKhhChDhEhF�hG�hKhHKubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubh�)��}�(h^NhKh>h�hDhEhG�h<�hh�h�hhAh�ubhj)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhihB�hKhhChDhEhF�hG�hKhHKubh)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAh�ubh�)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhb)��}�(h=KhKh>heh^NhDhEhF�hG�h<�h_KhhChAhfubhz)��}�(h^Nh<�h-K h=Kh_Kh>hvh@�hKhAh}hB�hKhhChDhEhF�hG�hHK ubhb)��}�(h=KhKh>heh^NhDhEhF�hG�h<�h_KhhChAhfubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhn)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAhqubh)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAh�ubhn)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAhqubh�)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubh7�Mace���)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubh�)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhj)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhihB�hKhhChDhEhF�hG�hKhHKubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubh7�Dagger���)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhO)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhNhB�hKhhChDhEhF�hG�hKhHKubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubh)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAh�ubhX�Cloth_Shirt���)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChA�Cloth Shirt�ubhj)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhihB�hKhhChDhEhF�hG�hKhHKubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubh)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAh�ubh�)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhs)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAhrhB�hKhhChDhEhF�hG�hKhHKubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhs)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAhrhB�hKhhChDhEhF�hG�hKhHKubh�)��}�(h=K#hKh>hehDhEhF�hG�h<�h_K#hhChAh�ubh��	Time_Bomb���)��}�(h<��radius�Kh>h<hK hA�Bomb��dur�KhKh�o�hDhE�damage�KhG��desc��Explodes up after 3 turns�ubhX�
Chain_Helm���)��}�(h=K
hKh>h]hDhEhF�hG�h<�h_KhhChA�
Chain Helm�ubh)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAh�ubh�)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubh)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAh�ubhZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ubh)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAh�ubh)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAh�ubh�)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubh7�Iron_Shield���)��}�(h^Nh<�h-K h=Kh_Kh>hvh@�hKhA�Iron Shield�hB�hKhhChDhEhF�hG�hHK ubh)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAh�ubh�)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhb)��}�(h=KhKh>heh^NhDhEhF�hG�h<�h_KhhChAhfubh�)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhn)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAhqubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhs)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAhrhB�hKhhChDhEhF�hG�hKhHKubh�)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhO)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhNhB�hKhhChDhEhF�hG�hKhHKubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubh�)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhj)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhihB�hKhhChDhEhF�hG�hKhHKubhj)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhihB�hKhhChDhEhF�hG�hKhHKubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubh)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAh�ubhj)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhihB�hKhhChDhEhF�hG�hKhHKubh�)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubh�)��}�(h^Nh<�h�Kh>h<hK hAh�h�KhKhh�hDhEj   KhG�j  j  ubh)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAh�ubh�)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubh�)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAh�ubh�)��}�(hKh>h�hDhEhG�h<�hh�h�hhAh�ubhz)��}�(h<�h-K h=Kh_Kh>hvh@�hKhAh}hB�hKhhChDhEhF�hG�hHK ubh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhn)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAhqubh�)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAh�ubh�)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubh�)��}�(h^NhKh>h�hDhEhG�h<�hh�h�hhAh�ubhb)��}�(h=KhKh>heh^NhDhEhF�hG�h<�h_KhhChAhfubhn)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAhqubhb)��}�(h=KhKh>heh^NhDhEhF�hG�h<�h_KhhChAhfubhs)��}�(h<�h-Kh=Kh>hvh@�hKhAhrhB�hKhhChDhEhF�hG�hKhHKubh�)��}�(h<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhj)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhihB�hKhhChDhEhF�hG�hKhHKubh��	GreenHerb���)��}�(h^Nh>h<hDhEhG�h<�h�+��healNum�KhA�
Green Herb�ubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhZ)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_K
hhChAh`ubhO)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhNhB�hKhhChDhEhF�hG�hKhHKubhb)��}�(h=KhKh>heh^NhDhEhF�hG�h<�h_KhhChAhfubhO)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhNhB�hKhhChDhEhF�hG�hKhHKubh�)��}�(h^Nh<�h�Kh>h<hK hAh�h�KhKhh�hDhEj   KhG�j  j  ubh�)��}�(h^Nh<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhn)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAhqubh�)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKube�exp�K��
baseHealth�M�
healthTemp�K �effects�]�h_K �	healthMax�M,�playerControlled���skillLevels�}�(hKhKhK h!Kh$K h'K h*K uhA�George�h^�Object�j�  ��)��}�(�col�KE�pLevel��LevelTypes.LevelTypes��Tower���)��}�(hh	�levelManager��LevelManager�j�  ��)��}�(�cursor�K �	levelList�]�j�  a�
messageSys��
MessageSys��Messages���)��}�(�retrieveLimit�K�messageLimit�M��messages�]�(�Goblin Grunt dropped Longsword��!Goblin Grunt dropped Leather Helm��Goblin Grunt dropped Buckler��!Goblin Grunt was killed by George��Goblin Grunt is afraid!��"George attacked Goblin Grunt for 4��Goblin Grunt missed George��George acquired 5 coins��"Goblin Grunt attacked George for 3��George picked up Bow�� Goblin Grunt picked up Cloth Hat�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 4��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George picked up Iron Helm��#Goblin Archer attacked George for 1��#Goblin Berserker dropped Gold Coins��&Goblin Berserker dropped Leather Shirt��"Goblin Berserker dropped Iron Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 4��#Goblin Archer attacked George for 1��&Goblin Berserker attacked George for 5��George acquired 12 coins��#Goblin Archer attacked George for 1��&Goblin Berserker attacked George for 5��George picked up Mace��#Goblin Archer attacked George for 1��$Goblin Berserker picked up Iron Helm��#Goblin Stonewall dropped Gold Coins��Goblin Stonewall dropped Mace��"Goblin Stonewall dropped Iron Helm��%Goblin Stonewall was killed by George��Goblin Stonewall is afraid!��&George attacked Goblin Stonewall for 2��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��&George attacked Goblin Berserker for 2��&George attacked Goblin Stonewall for 2��George used Fireball��&Goblin Stonewall attacked George for 3��&George attacked Goblin Berserker for 2��&George attacked Goblin Stonewall for 2��George used Lightning Bolt��George waited...��George waited...��George waited...��George picked up Bomb��George picked up Greatsword��George picked up Leather Shirt��George picked up Greatsword��George picked up Leather Helm��#Goblin Berserker dropped Greatsword��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 4��&Goblin Berserker attacked George for 5��&George attacked Goblin Berserker for 4��&Goblin Berserker attacked George for 5��George picked up Leather Helm��#Goblin Berserker dropped Greatsword��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 4��&Goblin Berserker attacked George for 5��George picked up Leather Helm��Goblin Berserker dropped Bomb��&Goblin Berserker dropped Leather Shirt��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 4��&Goblin Berserker attacked George for 5��George picked up Green Herb��&Goblin Berserker attacked George for 5��George picked up Spear��'Goblin Berserker picked up Leather Helm�� Goblin Lancer dropped Green Herb��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 4��Goblin Lancer missed George��#Goblin Lancer attacked George for 2��&George attacked Goblin Berserker for 2��&George attacked Goblin Berserker for 2��George used Fireball��#Goblin Lancer attacked George for 2��&George attacked Goblin Berserker for 2��#George attacked Goblin Lancer for 2��George used Lightning Bolt��George waited...��George waited...��George waited...��George acquired 8 coins��George picked up Bow��George acquired 8 coins��George picked up Longsword��George acquired 9 coins��George picked up Leather Shirt��George picked up Iron Helm��#Goblin Berserker dropped Gold Coins��&Goblin Berserker dropped Leather Shirt��"Goblin Berserker dropped Iron Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 4��&Goblin Berserker attacked George for 5��George acquired 5 coins��&Goblin Berserker attacked George for 5��George picked up Leather Shirt��$Goblin Berserker picked up Iron Helm��Goblin Grunt dropped Gold Coins��"Goblin Grunt dropped Leather Shirt��Goblin Grunt dropped Iron Helm��!Goblin Grunt was killed by George��Goblin Grunt is afraid!��"George attacked Goblin Grunt for 4��Goblin Grunt missed George��#George picked up Scroll of Fireball��"Goblin Grunt attacked George for 3��George picked up Mace�� Goblin Grunt picked up Iron Helm��+Goblin Stonewall dropped Scroll of Fireball��Goblin Stonewall dropped Mace��"Goblin Stonewall dropped Iron Helm��%Goblin Stonewall was killed by George��Goblin Stonewall is afraid!��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&George attacked Goblin Stonewall for 2��"George attacked Goblin Grunt for 2��George used Fireball��&George attacked Goblin Berserker for 2��George missed Goblin Grunt��&George attacked Goblin Stonewall for 2��George used Lightning Bolt��George acquired 8 coins��George picked up Cloth Shirt��George picked up Iron Helm��George picked up Dagger��George acquired 12 coins��George picked up Wooden Shield��#George picked up Scroll of Fireball��George picked up Cloth Shirt��George picked up Bow��George picked up Cloth Hat��George acquired 10 coins��George picked up Bomb��George acquired 13 coins��George acquired 12 coins��George picked up Bow��George picked up Spear��George picked up Cloth Hat��George picked up Leather Helm��George picked up Spear��George picked up Spear�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 6��George used Shocking Grasp��George used Shocking Grasp�� Goblin Lancer dropped Gold Coins��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 4��#Goblin Lancer attacked George for 2��George picked up Leather Helm��#Goblin Lancer attacked George for 2��#George attacked Goblin Lancer for 2��George used Lightning Bolt��#Goblin Lancer attacked George for 2��Goblin Lancer dropped Bomb��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 4��#Goblin Lancer attacked George for 2��#Goblin Lancer attacked George for 2��George picked up Leather Helm�� Goblin Lancer dropped Gold Coins��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 4��#Goblin Lancer attacked George for 2��#Goblin Archer attacked George for 1��#Goblin Lancer attacked George for 2��#Goblin Archer attacked George for 1��George waited...��#Goblin Archer attacked George for 1��George waited...��#Goblin Archer attacked George for 1��George waited...��#Goblin Archer attacked George for 1�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 4��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George waited...��George acquired 5 coins��George picked up Dagger��George picked up Leather Helm��Goblin Thief dropped Gold Coins��Goblin Thief dropped Dagger��!Goblin Thief dropped Leather Helm��!Goblin Thief was killed by George��"George attacked Goblin Thief for 2��George used Lightning Bolt��George used a Green Herb��George used a Green Herb��George used a Green Herb��George acquired 11 coins��George acquired 4 coins��George picked up Greatsword��George picked up Mace��George picked up Longsword��George picked up Leather Helm��Goblin Grunt dropped Gold Coins��Goblin Grunt dropped Longsword��!Goblin Grunt dropped Leather Helm��!Goblin Grunt was killed by George��Goblin Grunt is afraid!��"George attacked Goblin Grunt for 4��"Goblin Grunt attacked George for 3��George picked up Iron Helm��#Goblin Stonewall dropped Gold Coins��Goblin Stonewall dropped Mace��"Goblin Stonewall dropped Iron Helm��%Goblin Stonewall was killed by George��Goblin Stonewall is afraid!��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��Goblin Stonewall missed George��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&Goblin Stonewall attacked George for 3��George picked up Leather Helm��&George attacked Goblin Stonewall for 2��#Goblin Berserker dropped Greatsword��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 2��George used Fireball��&Goblin Berserker attacked George for 5��&George attacked Goblin Stonewall for 2��&George attacked Goblin Berserker for 2��George used Lightning Bolt��George waited...��"George attacked Goblin Grunt for 2��George used Lightning Bolt��"George attacked Goblin Thief for 2��&George attacked Goblin Berserker for 2��George used Fireball��George acquired 6 Arrows��George picked up Dagger��George picked up Leather Shirt��George picked up Bow��George picked up Cloth Hat��George picked up Iron Shield��Goblin Thief dropped Dagger��"Goblin Thief dropped Leather Shirt�� Goblin Thief dropped Iron Shield��!Goblin Thief was killed by George��"George attacked Goblin Thief for 2��George used Lightning Bolt��&Goblin Archer dropped Bundle of Arrows��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��#George attacked Goblin Archer for 2��"George attacked Goblin Thief for 2��George used Fireball��George acquired 14 coins��George picked up Bow��George picked up Cloth Hat�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��#George attacked Goblin Archer for 4��#Goblin Archer attacked George for 1��George acquired 10 coins��George picked up Cloth Hat��George picked up Leather Helm��George picked up Cloth Hat��George picked up Bow��George picked up Cloth Hat��"Goblin Thief picked up Iron Shield��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 4��George acquired 16 coins��George picked up Chain Helm��George picked up Bomb��George picked up Chain Shirt��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George picked up Longsword��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George picked up Leather Helm��#Goblin Archer attacked George for 1��Goblin Grunt dropped Longsword��!Goblin Grunt dropped Leather Helm��!Goblin Grunt was killed by George��Goblin Grunt is afraid!��"George attacked Goblin Grunt for 4��"George attacked Goblin Grunt for 2��George used Lightning Bolt��George waited...��George picked up Longsword��George acquired 12 coins��George picked up Bow��George picked up Cloth Hat�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 6��George used Shocking Grasp��George used Shocking Grasp��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George picked up Leather Helm��#Goblin Archer attacked George for 1��Goblin Archer is afraid!��#George attacked Goblin Archer for 2��Goblin Grunt dropped Longsword��!Goblin Grunt dropped Leather Helm��!Goblin Grunt was killed by George��Goblin Grunt is afraid!��"George attacked Goblin Grunt for 2��George used Fireball��Goblin Archer is afraid!��#George attacked Goblin Archer for 2��"George attacked Goblin Grunt for 2��George used Lightning Bolt��#Goblin Archer attacked George for 1��George waited...��#Goblin Archer attacked George for 1��George acquired 8 coins��George picked up Spear��George acquired 10 coins��George acquired 7 Arrows��George picked up Cloth Shirt��George picked up Cloth Hat��George picked up Leather Helm�� Goblin Lancer dropped Gold Coins��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 4��#Goblin Lancer attacked George for 2��#Goblin Lancer attacked George for 2��George waited...��#Goblin Lancer attacked George for 2��George picked up Greatsword��George picked up Leather Helm��#Goblin Berserker dropped Greatsword��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 6��George used Shocking Grasp��George used Shocking Grasp��George missed Goblin Lancer��George used Lightning Bolt��George acquired 5 coins��George picked up Dagger��George picked up Leather Helm��Goblin Thief dropped Gold Coins��Goblin Thief dropped Dagger��!Goblin Thief dropped Leather Helm��!Goblin Thief was killed by George��"George attacked Goblin Thief for 4��"Goblin Thief attacked George for 3��George waited...��George waited...��George waited...��George acquired 12 coins��George acquired 7 Arrows��George acquired 12 coins��George picked up Spear��George picked up Mace��George picked up Mace��George picked up Bow��George picked up Iron Helm��George leveled up!��)Goblin Stonewall dropped Bundle of Arrows��Goblin Stonewall dropped Mace��"Goblin Stonewall dropped Iron Helm��%Goblin Stonewall was killed by George��Goblin Stonewall is afraid!��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��Goblin Stonewall missed George��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��George picked up Cloth Hat��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 3��#Goblin Archer attacked George for 1��George picked up Iron Helm��#Goblin Stonewall dropped Gold Coins��Goblin Stonewall dropped Mace��"Goblin Stonewall dropped Iron Helm��%Goblin Stonewall was killed by George��Goblin Stonewall is afraid!��&George attacked Goblin Stonewall for 2��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��&George attacked Goblin Stonewall for 2��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��George missed Goblin Stonewall��#Goblin Archer attacked George for 1��&Goblin Stonewall attacked George for 3��George picked up Leather Helm�� Goblin Lancer dropped Gold Coins��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 3��#Goblin Lancer attacked George for 2��#George attacked Goblin Lancer for 3��#Goblin Lancer attacked George for 2��Goblin Lancer missed George��George acquired 7 coins��George picked up Leather Shirt��George picked up Wooden Shield��George acquired 5 coins��George picked up Leather Shirt��George picked up Bow��George picked up Cloth Hat�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 3��#Goblin Archer attacked George for 1��George picked up Spear��#Goblin Archer attacked George for 1��#Goblin Knight dropped Wooden Shield��#Goblin Knight dropped Leather Shirt��Goblin Knight dropped Spear��"Goblin Knight was killed by George��Goblin Knight is afraid!��#George attacked Goblin Knight for 3��#Goblin Knight attacked George for 4��#Goblin Archer attacked George for 1��#George attacked Goblin Knight for 3��#Goblin Knight attacked George for 4��#Goblin Archer attacked George for 1��George missed Goblin Knight��#Goblin Knight attacked George for 4��#Goblin Archer attacked George for 1��George missed Goblin Knight��Goblin Knight missed George��#Goblin Archer attacked George for 1��George missed Goblin Knight��#Goblin Knight attacked George for 4��#Goblin Archer attacked George for 1��#George picked up Scroll of Fireball��#Goblin Knight attacked George for 4��#Goblin Archer attacked George for 1��George picked up Leather Helm��#Goblin Knight attacked George for 4�� Goblin Archer dropped Gold Coins��#Goblin Archer dropped Leather Shirt��"Goblin Archer dropped Leather Helm��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 3��Goblin Knight picked up Spear��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George waited...��$Goblin Archer picked up Leather Helm��#Goblin Archer attacked George for 1��George picked up Greatsword��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George picked up Leather Helm��Goblin Archer missed George��#Goblin Archer attacked George for 1��#Goblin Berserker dropped Greatsword��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 3��#Goblin Archer attacked George for 1��&Goblin Berserker attacked George for 5��&George attacked Goblin Berserker for 3��#Goblin Archer attacked George for 1��&Goblin Berserker attacked George for 5��George missed Goblin Berserker��(Goblin Lancer dropped Scroll of Fireball��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 2��George used Lightning Bolt��&George attacked Goblin Berserker for 2��#George attacked Goblin Lancer for 2��George used Fireball��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George waited...��#Goblin Archer attacked George for 1��George acquired 11 coins��Goblin Archer missed George��George acquired 8 coins��George picked up Green Herb��George picked up Leather Shirt��George picked up Iron Helm��George acquired 11 coins��George picked up Greatsword��George waited...��George waited...��George acquired 8 coins��George picked up Leather Helm��#Goblin Berserker dropped Gold Coins��#Goblin Berserker dropped Greatsword��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 6��George used Shocking Grasp��George used Shocking Grasp��George picked up Leather Shirt��George picked up Leather Helm��#Goblin Berserker dropped Gold Coins��&Goblin Berserker dropped Leather Shirt��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 3��&Goblin Berserker attacked George for 5��George picked up Longsword��'Goblin Berserker picked up Leather Helm��George waited...��&George attacked Goblin Berserker for 2��Goblin Grunt dropped Longsword��!Goblin Grunt dropped Leather Helm��!Goblin Grunt was killed by George��Goblin Grunt is afraid!��"George attacked Goblin Grunt for 2��George used Fireball��"Goblin Grunt attacked George for 3��&George attacked Goblin Berserker for 2��"George attacked Goblin Grunt for 2��George used Lightning Bolt��George waited...��George waited...��George acquired 5 Arrows��George picked up Longsword��George acquired 6 coins��George acquired 4 coins��George picked up Bow��George picked up Bow��George picked up Cloth Hat�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 3��#Goblin Archer attacked George for 1��George picked up Cloth Hat��#Goblin Archer attacked George for 1�� Goblin Archer dropped Gold Coins��Goblin Archer dropped Bow��Goblin Archer dropped Cloth Hat��"Goblin Archer was killed by George��Goblin Archer is afraid!��#George attacked Goblin Archer for 3��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George missed Goblin Archer��Goblin Archer missed George��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��George picked up Iron Helm��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��&Goblin Knight dropped Bundle of Arrows��Goblin Knight dropped Longsword��Goblin Knight dropped Iron Helm��"Goblin Knight was killed by George��Goblin Knight is afraid!��#George attacked Goblin Knight for 3��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#Goblin Knight attacked George for 4��#George attacked Goblin Knight for 3��#Goblin Archer attacked George for 1��#Goblin Archer attacked George for 1��#George picked up Scroll of Fireball��George acquired 15 coins��George picked up Chain Shirt��George picked up Cloth Hat��George acquired 12 coins��George picked up Cloth Hat��George picked up Wooden Shield��George acquired 6 coins��George picked up Leather Shirt��George picked up Longsword��George picked up Iron Helm�� Goblin Knight dropped Gold Coins��Goblin Knight dropped Longsword��Goblin Knight dropped Iron Helm��"Goblin Knight was killed by George��Goblin Knight is afraid!��#George attacked Goblin Knight for 3��#Goblin Knight attacked George for 4��George picked up Spear��#Goblin Knight dropped Wooden Shield��#Goblin Knight dropped Leather Shirt��Goblin Knight dropped Spear��"Goblin Knight was killed by George��Goblin Knight is afraid!��#George attacked Goblin Knight for 3��#Goblin Knight attacked George for 4��#George attacked Goblin Knight for 3��#Goblin Knight attacked George for 4��George acquired 6 Arrows��#Goblin Knight attacked George for 4��George picked up Leather Shirt��Goblin Knight picked up Spear��)Goblin Berserker dropped Bundle of Arrows��&Goblin Berserker dropped Leather Shirt��Goblin Berserker dropped Spear��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 3��&Goblin Berserker attacked George for 5��George acquired 12 coins��&Goblin Berserker attacked George for 5��George picked up Leather Shirt��Goblin Berserker missed George��George picked up Leather Helm��&Goblin Berserker attacked George for 5��&George attacked Goblin Berserker for 2��#George attacked Goblin Knight for 2��#George attacked Goblin Knight for 2��George used Fireball��&Goblin Berserker attacked George for 5��George acquired 13 coins�� Goblin Berserker picked up Spear��George waited...��#Goblin Berserker dropped Gold Coins��&Goblin Berserker dropped Leather Shirt��%Goblin Berserker dropped Leather Helm��%Goblin Berserker was killed by George��Goblin Berserker is afraid!��&George attacked Goblin Berserker for 6��George used Shocking Grasp��George used Shocking Grasp��'Goblin Berserker picked up Leather Helm��&George attacked Goblin Berserker for 2��#George attacked Goblin Knight for 2��&George attacked Goblin Berserker for 2�� Goblin Lancer dropped Gold Coins��Goblin Lancer dropped Spear��"Goblin Lancer dropped Leather Helm��"Goblin Lancer was killed by George��Goblin Lancer is afraid!��#George attacked Goblin Lancer for 2��George used Lightning Bolt��#Goblin Lancer attacked George for 2��#Goblin Lancer attacked George for 2��George waited...��George waited...��#George attacked Goblin Lancer for 2��&George attacked Goblin Berserker for 2��George used Fireball��Player Ready: George��
Game Start�eub�	gameState�h�nextSeed�M7Bub�textWall��Cracked stone wall
��	textSpace��Dusty stone floor
��djikstra_Player_Away�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�h�     G�i      G�iP     G�i�     NNNNNNNNNNNNNNNNNG�k`     G�k�     G�k�     G�k�     G�l      G�lP     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK G�n      G�m�     G�m�     G�mp     G�m@     G�m     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�h�     G�h�     G�i      G�iP     NNNNNNNNNNNNNNNNNG�k0     G�k`     G�k�     G�k�     G�k�     G�l      NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�n      G�m�     G�m�     G�mp     G�m@     G�m     G�l�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�h0     G�h`     G�h�     G�h�     G�h�     G�i      NNNNNNNNNNNNNNNNNG�k      G�k0     G�k`     G�k�     G�k�     G�k�     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�m�     G�m�     G�mp     G�m@     G�m     G�l�     G�l�     G�l�     G�lP     G�l      G�k�     G�k�     G�k�     G�k`     G�k0     G�k      NNNNNNNNNNNNNNNNNNNG�i      G�h�     G�h�     G�h�     G�h`     G�h0     G�h      G�h0     G�h`     G�h�     G�h�     G�h�     NNNNNNNNNNNNNNNNNG�j�     G�k      G�k0     G�k`     G�k�     G�k�     G�k�     G�l      G�lP     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�n      G�m�     G�m�     G�mp     G�m@     G�m     G�l�     NNNNNNNNG�j�     NNNNNNNNNNNNNNNNNNNG�iP     NNNNNG�g�     G�h      G�h0     G�h`     G�h�     G�h�     NNNNNNNNNNNNNNNNNG�j�     G�j�     G�k      G�k0     G�k`     G�k�     G�k�     G�k�     G�l      NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK G�n      G�m�     G�m�     G�mp     G�m@     G�m     NNNNNNNNG�j�     NNNNNNNNNNNNNNNNNNNG�i�     NNNNNG�g�     G�g�     G�h      G�h0     G�h`     G�h�     G�h�     G�h�     G�i      G�iP     G�i�     G�i�     G�i�     G�j     G�j@     G�jp     NNNNNNNG�jp     G�j�     G�j�     G�k      G�k0     G�k`     G�k�     G�k�     G�k�     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�n      G�m�     G�m�     G�m�     G�m�     G�mp     G�m@     NNNNNNNNG�jp     NNNNG�i�     G�iP     G�i      G�h�     G�i      G�iP     NNNNNNNNNG�i�     NNNNNG�gp     NNNNNNNNNNNNNNG�j�     G�j�     G�k      G�k0     G�k      G�j�     G�j�     G�jp     G�j@     G�jp     G�j�     G�j�     G�k      G�k0     G�k`     G�k�     G�k�     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�m�     G�m�     G�mp     G�m�     G�m�     G�m�     G�mp     NNNNNNNNG�j@     G�j     G�i�     G�i�     G�i�     G�iP     G�i      G�h�     G�h�     G�h�     G�i      G�iP     G�i�     G�i�     G�i�     G�j     G�j@     G�jp     G�j@     G�j     G�i�     NNNNNG�g@     NNNNNNNNNNNNNNNNNNNNNNG�j     G�j@     G�jp     G�j�     G�j�     G�k      G�k0     G�k`     G�k�     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�m�     G�mp     G�m@     G�mp     G�m�     G�m�     G�m�     NNNNNNNNNNNNNG�i      G�h�     G�h�     G�h�     NNNNNNNNNNNNNNNNNG�g     NNNNNNNNNNNNNNNNNNNNNNG�i�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�mp     G�m@     G�m     G�m@     G�mp     G�m�     G�m�     NNNNNNNNNNNNNG�h�     G�h�     G�h�     G�h`     NNNNNNNNNNNNNNNNNG�f�     NNNNNNNNNNNNNNNNNNNNNNG�i�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�m@     G�m     G�l�     G�m     G�m@     G�mp     G�m�     NNNNNNNNNNNNNG�h�     G�h�     G�h`     G�h0     G�h`     G�h�     NNNNNNNNNNNNNNNG�f�     NNNNNNNNNNNNNNNNNNNNNNG�i�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�l�     NNNNNNNNNNNNNNNNNG�h�     G�h`     G�h0     G�h      G�h0     G�h`     NNNNNNNNNNNNNNNG�f�     NNNNNNNNNNNNNNNNNNNNNNG�iP     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�l�     NNNNNNNNNNNNNNNNNG�h`     G�h0     G�h      G�g�     G�h      G�h0     NNNNNNNNNNNNNNNG�fP     NNNNNNNNNNNNNNNNNNNNNNG�i      NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�lP     NNNNNNNNNNNNNNNNNG�h0     G�h      G�g�     G�g�     G�g�     G�h      NNNNNNNNNNNNNNNG�f      NNNNNNNNNNNNNNNNNNNNNNG�h�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�l      NNNNNNNNNNNNNNNNNNNNG�gp     NNNNNNNNNNNNNNNNNG�e�     G�e�     G�e�     G�e`     G�e0     G�e      G�d�     NNNNNNNNNNNNNNNNG�h�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�k�     NNNNNNNNNNNNNNNNNNNNG�g@     NNNNNNNNNNNNNNNNNNNNNNNG�d�     NNNNNNNNNNNNNNNNG�h�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�k�     NNNNNNNNNNNNNNNNNNNNG�g     NNNNNNNNNNNNNNNNNNNNNNNG�dp     NNNNNNNNNNNNNNNNG�h`     NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�k�     NNNNNNNNNNNNNNNNNNNNG�f�     G�f�     NNNNNNNNNNNNNNNNNNNNNNG�d@     NNNNNNNNNNNNNNNNG�h0     G�h      G�g�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�k`     NNNNNNNNNNNNNNNNNNNNNG�f�     NNNNNNNNNNNNNNNNNNNNNNG�d     NNNNNNNNNNNNNNNNNNG�g�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�j�     G�j�     G�k      G�k0     NNNNNNNNNNNNNNNNNNNNNG�fP     NNNNNNNNNNNNNNNNNNNNNNG�c�     NNNNNNNNNNNNNNNNNNG�gp     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�jp     NNNNNNNNNNNNNNNNNNG�e`     G�e0     G�e`     G�e�     G�e�     G�e�     G�f      G�fP     G�f�     G�f�     NNNNNNNNNNNNNNNNNNNG�c�     NNNNNNNNNNNNNNNNNNG�g@     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�j@     NNNNNNNNNNNNNNNNNNG�e0     G�e      G�e0     G�e`     G�e�     G�e�     G�e�     G�f      G�fP     G�f�     G�fP     G�f      G�e�     G�e�     G�e�     G�e`     G�e0     G�e      NNNNNNNNNNNG�c�     NNNNNNNNNNNNNNNNNNG�g     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�j     NNNNNNNNNNNNNNNNNNG�e      G�d�     G�e      G�e0     G�e`     G�e�     G�e�     G�e�     G�f      G�fP     NNNNNNNG�d�     NNNNNNNNNNNG�cP     NNNNNNNNNNNNNNNNNNG�f�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�j�     G�jp     G�j@     G�j     G�i�     G�i�     G�i�     G�iP     G�i�     NNNNNNNNNNNNNNG�d�     G�d�     G�d�     NNNNG�e�     G�e�     G�f      NNNNNNNG�d�     NNNNNNNNNNNG�c      NNNNNNNNNNNNNNNNG�fP     G�f�     G�f�     G�f�     G�f�     G�f�     G�g     G�g@     G�gp     G�g�     NNNNNNNNNNNNNNNNNNNe]�(NNG�jp     G�j@     G�j     G�i�     G�i�     G�i�     G�iP     G�i      G�iP     NNNNNNNNNNNNNNG�d�     G�dp     G�d�     NNNNG�e�     G�e�     G�e�     NNNNNNNG�dp     NNNNNNNNG�b�     G�b�     G�b�     G�b�     G�c      G�cP     G�c�     G�c�     G�c�     NNNNNNNNG�e�     G�e�     G�e�     G�f      G�fP     G�f�     G�f�     G�f�     G�f�     G�f�     G�g     G�g@     G�gp     NNNNNNNNNNNNNNNNNNNe]�(NNG�j@     G�j     G�i�     G�i�     G�i�     G�iP     G�i      G�h�     G�i      NNNNNNNNG�e�     G�e`     G�e0     G�e      G�d�     G�d�     G�dp     G�d@     G�dp     NNNNG�e`     G�e�     G�e�     NNNNNNNG�d@     NNNNNNNNG�b�     G�b`     G�b�     G�b�     G�b�     G�c      G�cP     G�c�     G�c�     NNNNNNNNG�e`     NNG�fP     G�f�     G�f�     G�f�     G�fP     G�f�     G�f�     G�f�     G�g     G�g@     NNNNNNNNNNNNNNNNNNNe]�(NNG�j     G�i�     G�i�     G�i�     G�iP     G�i      G�h�     G�h�     G�h�     NNNNNNNNG�e�     NNNNNG�d@     G�d     G�d@     NNNNG�e0     G�e`     G�e�     NNNNNNNG�d     G�c�     G�c�     G�c�     G�cP     G�c      G�b�     G�b�     G�b�     G�b`     G�b0     G�b`     G�b�     G�b�     G�b�     G�c      G�cP     G�c�     NNNNNNNNG�e0     NNG�f�     G�f�     G�f�     G�fP     G�f      G�fP     G�f�     G�f�     G�f�     G�g     NNNNNNNNNNNNNNNNNNNe]�(NNG�i�     G�i�     G�i�     G�iP     G�i      G�h�     G�h�     G�h�     G�h�     NNNNNNNNG�e�     NNNNNG�d     G�c�     G�d     G�d@     G�dp     G�d�     G�d�     G�e      G�e0     G�e`     NNNNNNNNNNNNNNNNG�b0     G�b      G�b0     G�b`     G�b�     G�b�     G�b�     G�c      G�cP     NNNNNNNNG�e      NNNNG�fP     G�f      G�e�     G�f      G�fP     G�f�     G�f�     G�f�     NNNNNNNNNNNNNNNNNNNe]�(NNG�j     G�i�     G�i�     NNNNG�h`     G�h�     NNNNNNNNG�f      NNNNNG�c�     G�c�     G�c�     G�d     G�d@     G�dp     G�d�     G�d�     G�e      G�e0     NNNNNNNNNNNNNNNNG�b      G�a�     G�b      G�b0     G�b`     G�b�     G�b�     G�b�     G�c      NNNNNNNNG�d�     NNNNG�f      G�e�     G�e�     G�e�     G�f      G�fP     G�f�     G�f�     NNNNNNNNNNNNNNNNNNNe]�(NNG�j@     G�j     G�i�     NNNNG�h0     G�h`     NNNNNNNNG�fP     NNNNNNG�c�     NNNNNNNNNNNNNNNNNNNNNNNNG�a�     G�a�     G�a�     G�b      G�b0     G�b`     G�b�     G�b�     G�b�     NNNNNNNNG�d�     NNNNNNG�e�     NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�jp     G�j@     G�j     NNNNG�h      G�h0     NNNNNNNNG�f�     NNNNNNG�cP     NNNNNNNNNNNNNNNNNNNNNNNNG�a�     G�ap     G�a�     G�a�     G�b      G�b0     G�b`     G�b�     G�b�     G�b�     G�c      G�cP     G�c�     G�c�     G�c�     G�d     G�d@     G�dp     NNNNNNG�e`     NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�j�     G�jp     G�j@     NNNNG�g�     G�h      G�h0     G�h      G�g�     G�g�     G�gp     G�g@     G�g     G�f�     G�f�     NNNNNNG�c      NNNNNNNNNNNNNNNNNNNNNNNNNG�a@     NNNNNNNNNNNNNNNNNNNNNNG�e0     G�e      G�d�     G�d�     G�dp     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�g�     NNNNNNNNNNNNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNNG�a     NNNNNNNNNNNNNNNNNNNNNNNNNNG�d@     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�gp     NNNNNNNNNNNNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNNG�`�     G�`�     G�`�     G�`P     G�`      NNNNNNNNNNNNNNNNNNNNNNG�d     NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�g@     NNNNNNNNNNNNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�_�     NNNNNNNNNNNNNNNNNNNNNNG�c�     NNNNNNNNNNNNNNNNNNNNe]�(NNNNG�f      G�fP     G�f�     G�f�     G�f�     G�g     NNNNNNNNNNNNNNNNG�b`     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�_�     NNNNNNNNNNNNNNNNNNNNNNG�c�     NNNNNNNNNNNNNNNNNNNNe]�(NNNNG�e�     NNNNNNNNNNNNNNNNNNNNNG�b0     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�_      NNNNNNNNNNNNNNNNNNNNNNG�c�     NNNNNNNNNNNNNNNNNNNNe]�(NNNNG�e�     NNNNNNNNNNNNNNNNNNNNNG�b      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�^�     NNNNNNNNNNNNNNNNNNNNG�cP     G�c�     G�cP     G�c      G�cP     NNNNNNNNNNNNNNNNNNe]�(NNNNG�e�     NNNNNNNNNNNNNNNNNNNNNG�a�     NNNNNNNNNNNNNNNNNNNNNNNG�_      G�^�     G�^`     G�^      G�]�     G�^      G�^`     G�^�     G�_      NNNNNNNNNNNNNNNNNNG�c      G�cP     G�c      G�b�     G�c      NNNNNNNNNNNNNNNNNNe]�(NNNNG�e`     NNNNNNNNNNNNNNNNNNNNNG�a�     NNNNNNNNNNNNNNNNNNNNNNNG�^�     G�^`     G�^      G�]�     G�]@     G�]�     G�^      G�^`     G�^�     NNNNNNNNNNNNNNNNNNG�b�     G�c      G�b�     G�b�     G�b�     NNNNNNNNNNNNNNNNNNe]�(NNNNG�e0     NNNNNNNNNNNNNNNNNNNNG�a�     G�ap     G�a@     G�a     G�a@     G�ap     G�a�     G�a�     G�b      NNNNNNNNNNNNNNNNG�^`     G�^      G�]�     G�]@     G�\�     G�]@     G�]�     G�^      G�^`     NNNNNNNNNNNNNNNG�b0     G�b`     G�b�     G�b�     G�b�     G�b�     G�b�     G�b�     NNNNNNNNNNNNNNNNNNe]�(NNNNG�e      NNNNNNNNNNNNNNG�b�     G�b`     G�b0     G�b      G�a�     G�a�     G�ap     G�a@     G�a     G�`�     G�a     G�a@     G�ap     G�a�     G�a�     NNNNNNNNNNNNNNNNG�^      G�]�     G�]@     G�\�     G�\�     G�\�     G�]@     G�]�     G�^      NNNNNNNNNNNNNNNG�b      G�b0     G�b`     G�b�     G�b�     G�b�     G�b`     G�b�     NNNNNNNNNNNNNNNNNNe]�(NNG�e0     G�e      G�d�     G�e      G�e0     G�e`     G�e�     G�e�     G�e�     NNNNNNNNG�b�     NNNNNG�a@     G�a     G�`�     G�`�     G�`�     G�a     G�a@     G�ap     G�a�     NNNNNNNNNNNNNNNNG�]�     G�]@     G�\�     G�\�     G�\      G�\�     G�\�     G�]@     G�]�     NNNNNNNNNG�`�     G�`�     G�a     G�a@     G�ap     G�a�     G�a�     G�b      G�b0     G�b`     G�b�     G�b`     G�b0     G�b`     NNNNNNNNNNNNNNNNNNe]�(NNG�e      G�d�     G�d�     G�d�     G�e      G�e0     G�e`     G�e�     G�e�     NNNNNNNNG�b�     NNNNNG�a     G�`�     G�`�     G�`�     G�`�     G�`�     G�a     G�a@     G�ap     NNNNNNNNNNNNNNNNG�]@     G�\�     G�\�     G�\      G�[�     G�\      G�\�     G�\�     G�]@     G�]�     G�^      G�^`     G�^�     G�_      G�_�     G�_�     G�`      G�`P     G�`�     NNNNNG�b      G�b0     G�b`     G�b�     G�b`     G�b0     G�b      G�b0     NNNNNNNNNNNNNNNNNNe]�(NNG�d�     G�d�     G�dp     G�d�     G�d�     G�e      G�e0     G�e`     G�e�     NNNNNNNNG�c      NNNNNG�`�     G�`�     G�`�     G�`P     G�`�     G�`�     G�`�     G�a     G�a@     NNNNNNNNNNNNNNNNG�\�     G�\�     G�\      G�[�     G�[`     G�[�     G�\      G�\�     G�\�     NNNNNNNNNNNNNNNG�b0     G�b`     G�b�     G�b`     G�b0     G�b      G�a�     G�b      NNNNNNNNNNNNNNNNNNe]�(NNG�d�     G�dp     G�d@     NNG�d�     G�e      G�e0     G�e`     NNNNNNNNG�cP     NNNNNG�`�     G�`�     G�`P     G�`      G�`P     G�`�     G�`�     G�`�     G�a     NNNNNNNNNNNNNNNNG�\�     G�\      G�[�     G�[`     G�[      G�[`     G�[�     G�\      G�\�     NNNNNNNNNNNNNNNNNNNNNG�a�     NNNNNNNNNNNNNNNNNNNe]�(NNG�dp     G�d@     G�d     NNG�d�     G�d�     G�e      G�e0     NNNNNNNNG�c�     NNNNNG�`�     G�`P     G�`      G�_�     G�`      G�`P     G�`�     G�`�     G�`�     NNNNNNNNNNNNNNNNG�\      G�[�     G�[`     G�[      G�Z�     G�[      G�[`     G�[�     G�\      NNNNNNNNNNNNNNNNNNNNNG�ap     NNNNNNNNNNNNNNNNNNNe]�(NNG�d@     G�d     G�c�     G�d     G�d@     G�dp     G�d�     G�d�     G�e      NNNNNNNNG�c�     NNNNNG�`P     G�`      G�_�     G�_�     G�_�     G�`      G�`P     G�`�     G�`�     NNNNNNNNNNNNNNNNG�[�     G�[`     G�[      G�Z�     G�Z@     G�Z�     G�[      G�[`     G�[�     NNNNNNNNNNNNNNNNNNNNNG�a@     NNNNNNNNNNNNNNNNNNNe]�(NNG�d     G�c�     G�c�     G�c�     G�d     G�d@     G�dp     G�d�     G�d�     NNNNNNNNG�c�     NNNNNG�`      G�_�     G�_�     G�_      G�_�     G�_�     G�`      G�`P     G�`�     NNNNNNNNNNNNNNNNNNNNG�Y�     NNNNNNNNNNNNNNNG�^`     G�^�     G�_      G�_�     G�_�     G�`      G�`P     G�`�     G�`�     G�`�     G�a     NNNNNNNNNNNNNNNNNNNe]�(NNG�c�     G�c�     G�c�     G�c�     G�c�     G�d     G�d@     G�dp     G�d�     G�d�     G�e      G�e0     G�e      G�d�     G�d�     G�dp     G�d@     G�d     NNNNNG�_�     G�_�     G�_      G�^�     G�_      G�_�     G�_�     G�`      G�`P     NNNNNNNNNNNNNNNNNNNNG�Y�     NNNNNNNNNNNNNNNG�^      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNG�cP     NNNNNNNNNNNNNNNNNNNNNNNG�^`     NNNNNNNNNNNNNNNNNNNNNNNNNG�Y      NNNNNNNNNNNNNNNG�]�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNG�c      G�b�     G�b�     G�b�     G�b`     NNNNNNNNNNNNNNNNNNNG�^      NNNNNNNNNNNNNNNNNNNNNNNNNG�X�     G�X`     G�X      G�W�     G�W@     NNNNNNNNNNNG�]@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNG�b0     NNNNNNNNNNNNNNNNNNNG�]�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�V�     NNNNNNNNNNNG�\�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNG�b      NNNNNNNNNNNNNNNNNNNG�]@     G�\�     G�\�     G�\      G�[�     NNNNNNNNNNNNNNNNNNNNNNNNNG�V�     NNNNNNNNNNNG�\�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�b�     G�b�     G�b�     G�b`     G�b0     G�b      G�a�     G�a�     G�ap     G�a@     NNNNNNNNNNNNNNNNNNNNG�[`     NNNNNNNNNNNNNNNNNNNNNNNNNG�V      NNNNNNNNNNNG�\      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�b�     G�b�     G�b`     G�b0     G�b      G�a�     G�a�     G�ap     G�a@     G�a     NNNNNNNNNNNNNNNNNNNNG�[      NNNNNNNNNNNNNNNNNNNNNNNNNG�U�     NNNNNNNNNNG�[`     G�[�     G�\      G�\�     G�\�     G�]@     G�]�     G�^      G�^`     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�b�     G�b`     G�b0     G�b      G�a�     G�a�     G�ap     G�a@     G�a     G�`�     G�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     NNNNNNNNNG�[      G�Z�     G�Z@     G�Z�     G�[      NNNNNNNNNNNNNNNNNNNNNNNNG�U`     NNNNNNNNNNG�[      G�[`     G�[�     G�\      G�\�     G�\�     G�]@     G�]�     G�^      NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�b�     G�b�     G�b`     G�b0     G�b      G�a�     G�a�     G�ap     G�a@     G�a     NNNNNNNG�^`     NNNNNNNNNG�Z�     G�Z@     G�Y�     G�Z@     G�Z�     NNNNNNNNNNNNNNNNNNG�S�     G�S      G�S�     G�S�     G�T@     G�T�     G�U      NNNNNNNNNNG�Z�     G�[      G�[`     G�[�     G�\      G�\�     G�\�     G�]@     G�]�     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�b�     G�b�     G�b�     G�b`     G�b0     G�b      NNNG�a@     NNNNNNNG�^      NNNNNNNG�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y�     G�Z@     NNNNNNNNNNNNNNNNNNG�S      G�R�     G�S      G�S�     G�S�     G�T@     G�T�     G�U      G�U`     G�U�     G�V      G�V�     G�V�     G�W@     G�W�     NNG�Z@     G�Z�     G�[      G�[`     G�[�     G�\      G�\�     G�\�     G�]@     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�c      G�b�     G�b�     G�b�     G�b`     G�b0     NNNG�ap     NNNNNNNG�]�     NNNNNNNG�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�Y�     G�Y�     NNNNNNNNNNNNNNNNNNG�R�     G�R`     G�R�     G�S      G�S�     G�S�     G�T@     NNNNNNNG�X      NNG�Y�     G�Z@     G�Z�     G�[      G�[`     G�[�     G�\      G�\�     G�\�     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�cP     G�c      G�b�     G�b�     G�b�     G�b`     NNNG�a�     NNNNNNNG�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�Y      G�Y�     NNNNNNNNNNNNNNNNNNG�R`     G�R      G�R`     G�R�     G�S      G�S�     G�S�     NNNNNNNG�X`     G�X�     G�Y      G�Y�     G�Y�     G�Z@     G�Z�     G�[      G�[`     G�[�     G�\      G�\�     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�c�     G�cP     G�c      G�b�     G�b�     G�b�     G�b`     G�b0     G�b      G�a�     NNNNNNNNNNNNNNNG�Y�     G�Y�     G�Y      G�X�     G�X`     G�X�     G�Y      NNNNNNNNNNNNNNNNNNG�R      G�Q�     G�R      G�R`     G�R�     G�S      G�S�     NNNNNNNNNNG�Y�     G�Z@     G�Z�     G�[      G�[`     G�[�     G�\      G�\�     G�\�     NNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNG�Y�     G�Y      G�X�     G�X`     G�X      G�X`     G�X�     NNNNNNNNNNNNNNNNNNG�Q�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�c      NNNNNNNNNNNNNNNNNNNNNNNNG�W�     NNNNNNNNNNNNNNNNNNNNG�Q@     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�cP     NNNNNNNNNNNNNNNNNNNNNNNNG�W@     NNNNNNNNNNNNNNNNNNNNG�P�     G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�c      NNNNNNNNNNNNNNNNNNNNNNNNG�V�     NNNNNNNNNNNNNNNNNNNNG�P�     G�P      G�P�     G�P�     G�Q@     G�Q�     G�R      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNG�V�     NNNNNNNNNNNNNNNNNNNNG�P      G�O�     G�P      G�P�     G�P�     G�Q@     G�Q�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�b0     G�b`     G�b�     G�b�     NNNNNNNNNNNNNNNNNNNNNNNNG�V      NNNNNNNNNNNNNNNNNNNNNG�N�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�b      NNNNNNNNNNNNNNNNNNNNNNNNNNNG�U�     NNNNNNNNNNNNNNNNNNNNNG�N      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�a�     NNNNNNNNNNNNNNNNNNNNNNNNNG�T�     G�U      G�U`     NNNNNNNNNNNNNNNNNNNNNG�M@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�a�     NNNNNNNNNNNNNNNNNNNNNNNNNG�T@     NNNNNNNNNNNNNNNNNNNNNNNG�L�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�ap     NNNNNNNNNNNNNNNNNNNNNNNNNG�S�     NNNNNNNNNNNNNNNNNG�G@     G�H      G�H�     G�I�     G�J@     G�K      G�K�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�a@     NNNNNNNNNNNNNNNNNNNNNG�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     NNNNNNNNNNNNNNG�F�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�a@     G�a     G�`�     G�`�     G�`�     G�`P     G�`      NNNNNNNNNNNNNNNNG�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      NNNNNNNNNG�E�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�a     G�`�     G�`�     G�`�     G�`P     G�`      G�_�     NNNNNNNNNNNNNNNNG�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     NNNNG�O�     NNNNNNNNNG�E      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`�     G�`�     G�`P     G�`      G�_�     G�_�     NNNNNNNNNNNNNNNNG�U`     G�U      NNNG�S�     G�S      G�R�     NNNNG�N�     NNNNNNNNNG�D@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      NNNNNNNNNNNNNNNNG�U�     G�U`     NNNG�S�     G�S�     G�S      NNNNG�N      NNNNNNNNG�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     NNNNNNNNNNNNNNNNG�V      G�U�     NNNG�T@     G�S�     G�S�     NNNNG�M@     NNNNNNNNG�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     NNNNNNNNNNNNNNNNNG�      G�"      G�%      G�(      G�+      G�.      G�0�     G�2      G�3�     G�5      NNNNNNNNNNNNNNNNNNNe]�(NNG�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     NNNNNNNNG�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     NNNNG�L�     NNNNNNNNG�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      NNNNNNNNNNNNNNNNNG�      G�      G�"      G�%      G�(      G�+      G�.      G�0�     G�2      G�3�     NNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`P     NNG�^�     G�^`     G�^      NNNNNNNNG�Y�     NNNNNNNG�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     NNNNG�K�     NNNNNNNNG�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�(      G�%      G�"      NNNNNNG�      G�      G�      G�"      G�%      G�(      G�+      G�.      G�0�     G�2      NNNNNNNNNNNNNNNNNNNe]�(NNG�`P     G�`      NNG�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     NNNNNNNNNNNNNNNNNNNG�K      NNNNNNNNG�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      NNNNNNNNNNG�      G�      G�      G�      G��      G�       G��      G�      G�      G�      G�      G�"      G�%      G�(      G�+      G�.      G�0�     NNNNNNNNNNNNNNNNNNNe]�(NNG�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      NNNNNNNNNNNNNNNNNNNNNNNNNNNNG�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     NNNNNNNNNNNNNNNNNG�      G�      G�      G�"      G�%      G�(      G�+      G�.      G�0�     G�2      NNNNNNNNNNNNNNNNNNNe]�(NNG�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�B      G�A@     G�@�     G�?�     G�>      NNNNNNNNNNNNNNNNNG�      G�      G�"      G�%      G�(      G�+      G�.      G�0�     G�2      G�3�     NNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�B�     G�B      G�A@     G�@�     G�?�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�C�     G�B�     G�B      G�A@     G�@�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�consumeList�]�(jf  h��Bundle_Of_Arrows���h��
Gold_Coins���h�h�e�Tiles�}�(K }�(K �Tile�j  ��)��}�(j�  K �Objects�]�j�  j�  �row�K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubK j  )��}�(j�  K j  ]�j�  j�  j  K ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K ubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  �      ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�KGaj�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�Kaj�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�Kaj�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK	}�(K j  )��}�(j�  K j  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K	ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubKj  )��}�(j�  Kj  ]�j�  j�  j  K	ubK j  )��}�(j�  K j  ]�j�  j�  j  K	ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K	ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K	ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K	ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K	ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K	ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K	ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K	ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K	ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K	ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K	ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K	ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K	ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K	ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K	ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K	ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K	ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K	ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K	ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K	ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K	ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K	ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K	ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K	ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K	ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K	ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K	ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K	ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K	ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K	ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K	ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K	ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K	ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K	ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K	ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K	ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K	ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K	ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K	ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K	ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K	ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K	ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K	ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K	ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K	ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K	ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K	ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K	ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K	ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K	ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K	ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K	ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K	ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K	ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K	ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K	ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K	ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K	ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K	ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K	ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K	ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K	ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K	ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K	ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K	ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K	ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K	ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K	ubuK
}�(K j  )��}�(j�  K j  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K
ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubKj  )��}�(j�  Kj  ]�j�  j�  j  K
ubK j  )��}�(j�  K j  ]�j�  j�  j  K
ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K
ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K
ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K
ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K
ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K
ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K
ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K
ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K
ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K
ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K
ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K
ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K
ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K
ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K
ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K
ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K
ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K
ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K
ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K
ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K
ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K
ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K
ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K
ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K
ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K
ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K
ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K
ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K
ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K
ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K
ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K
ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K
ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K
ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K
ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K
ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K
ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K
ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K
ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K
ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K
ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K
ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K
ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K
ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K
ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K
ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K
ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K
ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K
ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K
ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K
ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K
ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K
ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K
ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K
ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K
ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K
ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K
ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K
ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K
ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K
ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K
ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K
ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K
ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K
ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K
ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K
ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K
ubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�Kaj�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�Kaj�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  �      )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  �      KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK	j  )��}�(j�  K	j  ]�j�  j�  j  KubK
j  )��}�(j�  K
j  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubKj  )��}�(j�  Kj  ]�j�  j�  j  KubK j  )��}�(j�  K j  ]�j�  j�  j  KubK!j  )��}�(j�  K!j  ]�j�  j�  j  KubK"j  )��}�(j�  K"j  ]�j�  j�  j  KubK#j  )��}�(j�  K#j  ]�j�  j�  j  KubK$j  )��}�(j�  K$j  ]�j�  j�  j  KubK%j  )��}�(j�  K%j  ]�j�  j�  j  KubK&j  )��}�(j�  K&j  ]�j�  j�  j  KubK'j  )��}�(j�  K'j  ]�j�  j�  j  KubK(j  )��}�(j�  K(j  ]�j�  j�  j  KubK)j  )��}�(j�  K)j  ]�j�  j�  j  KubK*j  )��}�(j�  K*j  ]�j�  j�  j  KubK+j  )��}�(j�  K+j  ]�j�  j�  j  KubK,j  )��}�(j�  K,j  ]�j�  j�  j  KubK-j  )��}�(j�  K-j  ]�j�  j�  j  KubK.j  )��}�(j�  K.j  ]�j�  j�  j  KubK/j  )��}�(j�  K/j  ]�j�  j�  j  KubK0j  )��}�(j�  K0j  ]�j�  j�  j  KubK1j  )��}�(j�  K1j  ]�j�  j�  j  KubK2j  )��}�(j�  K2j  ]�j�  j�  j  KubK3j  )��}�(j�  K3j  ]�j�  j�  j  KubK4j  )��}�(j�  K4j  ]�j�  j�  j  KubK5j  )��}�(j�  K5j  ]�j�  j�  j  KubK6j  )��}�(j�  K6j  ]�j�  j�  j  KubK7j  )��}�(j�  K7j  ]�j�  j�  j  KubK8j  )��}�(j�  K8j  ]�j�  j�  j  KubK9j  )��}�(j�  K9j  ]�j�  j�  j  KubK:j  )��}�(j�  K:j  ]�j�  j�  j  KubK;j  )��}�(j�  K;j  ]�j�  j�  j  KubK<j  )��}�(j�  K<j  ]�j�  j�  j  KubK=j  )��}�(j�  K=j  ]�j�  j�  j  KubK>j  )��}�(j�  K>j  ]�j�  j�  j  KubK?j  )��}�(j�  K?j  ]�j�  j�  j  KubK@j  )��}�(j�  K@j  ]�j�  j�  j  KubKAj  )��}�(j�  KAj  ]�j�  j�  j  KubKBj  )��}�(j�  KBj  ]�j�  j�  j  KubKCj  )��}�(j�  KCj  ]�j�  j�  j  KubKDj  )��}�(j�  KDj  ]�j�  j�  j  KubKEj  )��}�(j�  KEj  ]�j�  j�  j  KubKFj  )��}�(j�  KFj  ]�j�  j�  j  KubKGj  )��}�(j�  KGj  ]�j�  j�  j  KubKHj  )��}�(j�  KHj  ]�j�  j�  j  KubKIj  )��}�(j�  KIj  ]�j�  j�  j  KubKJj  )��}�(j�  KJj  ]�j�  j�  j  KubKKj  )��}�(j�  KKj  ]�j�  j�  j  KubKLj  )��}�(j�  KLj  ]�j�  j�  j  KubKMj  )��}�(j�  KMj  ]�j�  j�  j  KubKNj  )��}�(j�  KNj  ]�j�  j�  j  KubKOj  )��}�(j�  KOj  ]�j�  j�  j  KubKPj  )��}�(j�  KPj  ]�j�  j�  j  KubKQj  )��}�(j�  KQj  ]�j�  j�  j  KubKRj  )��}�(j�  KRj  ]�j�  j�  j  KubKSj  )��}�(j�  KSj  ]�j�  j�  j  KubKTj  )��}�(j�  KTj  ]�j�  j�  j  KubKUj  )��}�(j�  KUj  ]�j�  j�  j  KubKVj  )��}�(j�  KVj  ]�j�  j�  j  KubKWj  )��}�(j�  KWj  ]�j�  j�  j  KubKXj  )��}�(j�  KXj  ]�j�  j�  j  KubKYj  )��}�(j�  KYj  ]�j�  j�  j  KubKZj  )��}�(j�  KZj  ]�j�  j�  j  KubK[j  )��}�(j�  K[j  ]�j�  j�  j  KubK\j  )��}�(j�  K\j  ]�j�  j�  j  KubK]j  )��}�(j�  K]j  ]�j�  j�  j  KubK^j  )��}�(j�  K^j  ]�j�  j�  j  KubK_j  )��}�(j�  K_j  ]�j�  j�  j  KubK`j  )��}�(j�  K`j  ]�j�  j�  j  KubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KubuK }�(K j  )��}�(j�  K j  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubKj  )��}�(j�  Kj  ]�j�  j�  j  K ubK j  )��}�(j�  K j  ]�j�  j�  j  K ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K ubuK!}�(K j  )��}�(j�  K j  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K!ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubKj  )��}�(j�  Kj  ]�j�  j�  j  K!ubK j  )��}�(j�  K j  ]�j�  j�  j  K!ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K!ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K!ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K!ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K!ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K!ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K!ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K!ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K!ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K!ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K!ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K!ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K!ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K!ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K!ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K!ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K!ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K!ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K!ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K!ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K!ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K!ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K!ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K!ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K!ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K!ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K!ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K!ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K!ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K!ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K!ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K!ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K!ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K!ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K!ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K!ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K!ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K!ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K!ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K!ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K!ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K!ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K!ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K!ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K!ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K!ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K!ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K!ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K!ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K!ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K!ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K!ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K!ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K!ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K!ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K!ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K!ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K!ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K!ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K!ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K!ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K!ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K!ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K!ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K!ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K!ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K!ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K!ubuK"}�(K j  )��}�(j�  K j  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K"ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubKj  )��}�(j�  Kj  ]�j�  j�  j  K"ubK j  )��}�(j�  K j  ]�j�  j�  j  K"ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K"ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K"ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K"ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K"ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K"ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K"ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K"ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K"ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K"ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K"ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K"ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K"ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K"ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K"ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K"ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K"ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K"ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K"ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K"ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K"ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K"ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K"ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K"ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K"ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K"ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K"ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K"ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K"ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K"ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K"ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K"ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K"ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K"ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K"ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K"ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K"ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K"ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K"ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K"ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K"ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K"ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K"ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K"ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K"ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K"ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K"ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K"ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K"ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K"ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K"ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K"ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K"ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K"ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K"ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K"ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K"ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K"ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K"ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K"ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K"ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K"ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K"ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K"ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K"ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K"ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K"ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K"ubuK#}�(K j  )��}�(j�  K j  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K#ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubKj  )��}�(j�  Kj  ]�j�  j�  j  K#ubK j  )��}�(j�  K j  ]�j�  j�  j  K#ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K#ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K#ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K#ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K#ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K#ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K#ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K#ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K#ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K#ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K#ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K#ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K#ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K#ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K#ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K#ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K#ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K#ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K#ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K#ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K#ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K#ubK6j  )��}�(j�  K6j  ]�K#aj�  j�  j  K#ubK7j  )��}�(j�  K7j  ]�K$aj�  j�  j  K#ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K#ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K#ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K#ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K#ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K#ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K#ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K#ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K#ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K#ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K#ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K#ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K#ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K#ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K#ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K#ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K#ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K#ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K#ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K#ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K#ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K#ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K#ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K#ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K#ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K#ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K#ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K#ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K#ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K#ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K#ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K#ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K#ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K#ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K#ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K#ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K#ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K#ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K#ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K#ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K#ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K#ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K#ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K#ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K#ubuK$}�(K j  )��}�(j�  K j  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K$ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubKj  )��}�(j�  Kj  ]�j�  j�  j  K$ubK j  )��}�(j�  K j  ]�j�  j�  j  K$ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K$ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K$ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K$ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K$ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K$ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K$ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K$ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K$ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K$ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K$ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K$ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K$ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K$ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K$ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K$ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K$ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K$ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K$ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K$ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K$ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K$ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K$ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K$ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K$ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K$ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K$ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K$ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K$ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K$ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K$ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K$ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K$ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K$ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K$ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K$ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K$ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K$ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K$ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K$ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K$ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K$ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K$ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K$ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K$ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K$ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K$ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K$ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K$ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K$ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K$ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K$ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K$ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K$ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K$ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K$ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K$ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K$ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K$ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K$ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K$ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K$ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K$ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K$ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K$ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K$ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K$ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K$ubuK%}�(K j  )��}�(j�  K j  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K%ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubKj  )��}�(j�  Kj  ]�j�  j�  j  K%ubK j  )��}�(j�  K j  ]�j�  j�  j  K%ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K%ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K%ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K%ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K%ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K%ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K%ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K%ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K%ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K%ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K%ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K%ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K%ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K%ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K%ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K%ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K%ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K%ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K%ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K%ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K%ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K%ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K%ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K%ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K%ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K%ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K%ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K%ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K%ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K%ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K%ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K%ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K%ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K%ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K%ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K%ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K%ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K%ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K%ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K%ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K%ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K%ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K%ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K%ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K%ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K%ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K%ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K%ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K%ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K%ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K%ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K%ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K%ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K%ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K%ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K%ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K%ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K%ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K%ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K%ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K%ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K%ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K%ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K%ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K%ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K%ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K%ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K%ubuK&}�(K j  )��}�(j�  K j  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K&ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubKj  )��}�(j�  Kj  ]�j�  j�  j  K&ubK j  )��}�(j�  K j  ]�j�  j�  j  K&ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K&ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K&ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K&ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K&ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K&ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K&ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K&ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K&ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K&ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K&ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K&ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K&ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K&ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K&ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K&ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K&ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K&ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K&ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K&ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K&ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K&ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K&ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K&ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K&ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K&ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K&ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K&ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K&ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K&ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K&ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K&ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K&ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K&ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K&ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K&ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K&ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K&ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K&ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K&ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K&ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K&ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K&ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K&ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K&ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K&ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K&ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K&ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K&ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K&ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K&ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K&ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K&ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K&ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K&ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K&ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K&ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K&ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K&ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K&ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K&ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K&ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K&ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K&ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K&ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K&ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K&ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K&ubuK'}�(K j  )��}�(j�  K j  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K'ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubKj  )��}�(j�  Kj  ]�j�  j�  j  K'ubK j  )��}�(j�  K j  ]�j�  j�  j  K'ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K'ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K'ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K'ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K'ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K'ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K'ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K'ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K'ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K'ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K'ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K'ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K'ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K'ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K'ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K'ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K'ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K'ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K'ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K'ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K'ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K'ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K'ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K'ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K'ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K'ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K'ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K'ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K'ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K'ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K'ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K'ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K'ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K'ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K'ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K'ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K'ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K'ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K'ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K'ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K'ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K'ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K'ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K'ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K'ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K'ubKNj  )��}�(j�  KNj  ]�K�aj�  j�  j  K'ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K'ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K'ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K'ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K'ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K'ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K'ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K'ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K'ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K'ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K'ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K'ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K'ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K'ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K'ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K'ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K'ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K'ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K'ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K'ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K'ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K'ubuK(}�(K j  )��}�(j�  K j  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K(ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubKj  )��}�(j�  Kj  ]�j�  j�  j  K(ubK j  )��}�(j�  K j  ]�j�  j�  j  K(ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K(ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K(ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K(ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K(ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K(ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K(ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K(ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K(ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K(ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K(ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K(ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K(ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K(ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K(ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K(ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K(ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K(ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K(ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K(ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K(ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K(ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K(ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K(ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K(ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K(ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K(ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K(ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K(ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K(ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K(ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K(ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K(ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K(ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K(ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K(ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K(ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K(ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K(ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K(ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K(ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K(ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K(ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K(ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K(ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K(ubKNj  )��}�(j�  KNj  ]�K'aj�  j�  j  K(ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K(ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K(ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K(ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K(ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K(ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K(ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K(ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K(ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K(ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K(ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K(ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K(ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K(ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K(ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K(ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K(ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K(ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K(ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K(ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K(ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K(ubuK)}�(K j  )��}�(j�  K j  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K)ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubKj  )��}�(j�  Kj  ]�j�  j�  j  K)ubK j  )��}�(j�  K j  ]�j�  j�  j  K)ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K)ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K)ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K)ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K)ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K)ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K)ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K)ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K)ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K)ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K)ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K)ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K)ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K)ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K)ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K)ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K)ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K)ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K)ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K)ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K)ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K)ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K)ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K)ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K)ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K)ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K)ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K)ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K)ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K)ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K)ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K)ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K)ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K)ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K)ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K)ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K)ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K)ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K)ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K)ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K)ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K)ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K)ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K)ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K)ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K)ubKNj  )��}�(j�  KNj  ]�K*aj�  j�  j  K)ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K)ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K)ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K)ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K)ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K)ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K)ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K)ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K)ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K)ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K)ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K)ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K)ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K)ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K)ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K)ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K)ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K)ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K)ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K)ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K)ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K)ubuK*}�(K j  )��}�(j�  K j  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K*ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubKj  )��}�(j�  Kj  ]�j�  j�  j  K*ubK j  )��}�(j�  K j  ]�j�  j�  j  K*ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K*ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K*ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K*ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K*ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K*ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K*ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K*ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K*ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K*ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K*ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K*ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K*ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K*ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K*ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K*ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K*ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K*ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K*ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K*ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K*ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K*ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K*ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K*ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K*ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K*ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K*ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K*ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K*ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K*ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K*ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K*ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K*ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K*ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K*ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K*ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K*ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K*ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K*ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K*ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K*ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K*ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K*ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K*ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K*ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K*ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K*ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K*ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K*ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K*ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K*ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K*ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K*ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K*ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K*ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K*ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K*ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K*ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K*ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K*ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K*ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K*ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K*ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K*ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K*ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K*ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K*ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K*ubuK+}�(K j  )��}�(j�  K j  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K+ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubKj  )��}�(j�  Kj  ]�j�  j�  j  K+ubK j  )��}�(j�  K j  ]�j�  j�  j  K+ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K+ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K+ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K+ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K+ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K+ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K+ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K+ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K+ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K+ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K+ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K+ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K+ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K+ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K+ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K+ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K+ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K+ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K+ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K+ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K+ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K+ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K+ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K+ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K+ubK9j  )��}�(j�  K9j  ]�K,aj�  j�  j  K+ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K+ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K+ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K+ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K+ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K+ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K+ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K+ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K+ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K+ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K+ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K+ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K+ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K+ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K+ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K+ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K+ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K+ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K+ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K+ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K+ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K+ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K+ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K+ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K+ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K+ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K+ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K+ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K+ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K+ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K+ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K+ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K+ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K+ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K+ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K+ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K+ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K+ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K+ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K+ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K+ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K+ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K+ubuK,}�(K j  )��}�(j�  K j  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�K/aj�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�K0aj�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K,ubK
j  )��}�(j�  K
j  ]�K1aj�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )��}�(j�  Kj  ]�j�  j�  j  K,ubKj  )���      }�(j�  Kj  ]�j�  j�  j  K,ubK j  )��}�(j�  K j  ]�j�  j�  j  K,ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K,ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K,ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K,ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K,ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K,ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K,ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K,ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K,ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K,ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K,ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K,ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K,ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K,ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K,ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K,ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K,ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K,ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K,ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K,ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K,ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K,ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K,ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K,ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K,ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K,ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K,ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K,ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K,ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K,ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K,ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K,ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K,ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K,ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K,ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K,ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K,ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K,ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K,ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K,ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K,ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K,ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K,ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K,ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K,ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K,ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K,ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K,ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K,ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K,ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K,ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K,ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K,ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K,ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K,ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K,ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K,ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K,ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K,ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K,ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K,ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K,ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K,ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K,ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K,ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K,ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K,ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K,ubuK-}�(K j  )��}�(j�  K j  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K-ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�K3aj�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubKj  )��}�(j�  Kj  ]�j�  j�  j  K-ubK j  )��}�(j�  K j  ]�j�  j�  j  K-ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K-ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K-ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K-ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K-ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K-ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K-ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K-ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K-ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K-ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K-ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K-ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K-ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K-ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K-ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K-ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K-ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K-ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K-ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K-ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K-ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K-ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K-ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K-ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K-ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K-ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K-ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K-ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K-ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K-ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K-ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K-ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K-ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K-ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K-ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K-ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K-ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K-ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K-ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K-ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K-ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K-ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K-ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K-ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K-ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K-ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K-ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K-ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K-ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K-ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K-ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K-ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K-ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K-ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K-ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K-ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K-ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K-ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K-ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K-ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K-ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K-ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K-ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K-ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K-ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K-ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K-ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K-ubuK.}�(K j  )��}�(j�  K j  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K.ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubKj  )��}�(j�  Kj  ]�j�  j�  j  K.ubK j  )��}�(j�  K j  ]�j�  j�  j  K.ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K.ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K.ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K.ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K.ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K.ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K.ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K.ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K.ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K.ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K.ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K.ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K.ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K.ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K.ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K.ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K.ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K.ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K.ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K.ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K.ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K.ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K.ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K.ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K.ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K.ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K.ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K.ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K.ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K.ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K.ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K.ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K.ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K.ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K.ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K.ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K.ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K.ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K.ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K.ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K.ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K.ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K.ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K.ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K.ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K.ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K.ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K.ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K.ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K.ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K.ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K.ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K.ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K.ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K.ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K.ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K.ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K.ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K.ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K.ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K.ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K.ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K.ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K.ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K.ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K.ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K.ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K.ubuK/}�(K j  )��}�(j�  K j  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�K8aj�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K/ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubKj  )��}�(j�  Kj  ]�j�  j�  j  K/ubK j  )��}�(j�  K j  ]�j�  j�  j  K/ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K/ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K/ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K/ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K/ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K/ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K/ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K/ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K/ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K/ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K/ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K/ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K/ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K/ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K/ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K/ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K/ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K/ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K/ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K/ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K/ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K/ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K/ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K/ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K/ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K/ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K/ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K/ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K/ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K/ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K/ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K/ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K/ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K/ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K/ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K/ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K/ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K/ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K/ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K/ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K/ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K/ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K/ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K/ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K/ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K/ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K/ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K/ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K/ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K/ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K/ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K/ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K/ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K/ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K/ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K/ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K/ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K/ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K/ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K/ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K/ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K/ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K/ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K/ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K/ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K/ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K/ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K/ubuK0}�(K j  )��}�(j�  K j  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K0ubK
j  )��}�(j�  K
j  ]�K:aj�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubKj  )��}�(j�  Kj  ]�j�  j�  j  K0ubK j  )��}�(j�  K j  ]�j�  j�  j  K0ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K0ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K0ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K0ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K0ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K0ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K0ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K0ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K0ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K0ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K0ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K0ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K0ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K0ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K0ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K0ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K0ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K0ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K0ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K0ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K0ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K0ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K0ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K0ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K0ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K0ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K0ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K0ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K0ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K0ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K0ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K0ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K0ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K0ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K0ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K0ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K0ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K0ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K0ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K0ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K0ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K0ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K0ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K0ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K0ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K0ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K0ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K0ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K0ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K0ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K0ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K0ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K0ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K0ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K0ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K0ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K0ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K0ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K0ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K0ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K0ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K0ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K0ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K0ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K0ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K0ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K0ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K0ubuK1}�(K j  )��}�(j�  K j  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K1ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�K=aj�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubKj  )��}�(j�  Kj  ]�j�  j�  j  K1ubK j  )��}�(j�  K j  ]�j�  j�  j  K1ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K1ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K1ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K1ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K1ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K1ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K1ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K1ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K1ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K1ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K1ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K1ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K1ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K1ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K1ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K1ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K1ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K1ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K1ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K1ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K1ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K1ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K1ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K1ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K1ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K1ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K1ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K1ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K1ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K1ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K1ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K1ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K1ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K1ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K1ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K1ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K1ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K1ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K1ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K1ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K1ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K1ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K1ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K1ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K1ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K1ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K1ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K1ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K1ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K1ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K1ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K1ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K1ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K1ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K1ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K1ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K1ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K1ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K1ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K1ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K1ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K1ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K1ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K1ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K1ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K1ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K1ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K1ubuK2}�(K j  )��}�(j�  K j  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K2ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubKj  )��}�(j�  Kj  ]�j�  j�  j  K2ubK j  )��}�(j�  K j  ]�j�  j�  j  K2ubK!j  )��}�(j�  K!j  ]�K>aj�  j�  j  K2ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K2ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K2ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K2ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K2ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K2ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K2ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K2ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K2ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K2ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K2ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K2ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K2ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K2ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K2ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K2ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K2ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K2ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K2ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K2ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K2ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K2ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K2ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K2ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K2ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K2ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K2ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K2ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K2ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K2ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K2ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K2ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K2ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K2ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K2ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K2ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K2ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K2ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K2ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K2ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K2ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K2ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K2ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K2ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K2ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K2ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K2ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K2ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K2ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K2ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K2ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K2ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K2ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K2ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K2ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K2ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K2ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K2ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K2ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K2ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K2ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K2ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K2ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K2ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K2ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K2ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K2ubuK3}�(K j  )��}�(j�  K j  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K3ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubKj  )��}�(j�  Kj  ]�j�  j�  j  K3ubK j  )��}�(j�  K j  ]�j�  j�  j  K3ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K3ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K3ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K3ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K3ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K3ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K3ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K3ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K3ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K3ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K3ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K3ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K3ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K3ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K3ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K3ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K3ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K3ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K3ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K3ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K3ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K3ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K3ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K3ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K3ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K3ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K3ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K3ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K3ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K3ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K3ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K3ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K3ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K3ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K3ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K3ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K3ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K3ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K3ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K3ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K3ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K3ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K3ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K3ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K3ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K3ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K3ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K3ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K3ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K3ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K3ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K3ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K3ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K3ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K3ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K3ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K3ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K3ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K3ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K3ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K3ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K3ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K3ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K3ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K3ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K3ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K3ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K3ubuK4}�(K j  )��}�(j�  K j  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K4ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubKj  )��}�(j�  Kj  ]�j�  j�  j  K4ubK j  )��}�(j�  K j  ]�j�  j�  j  K4ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K4ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K4ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K4ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K4ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K4ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K4ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K4ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K4ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K4ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K4ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K4ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K4ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K4ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K4ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K4ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K4ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K4ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K4ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K4ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K4ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K4ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K4ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K4ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K4ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K4ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K4ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K4ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K4ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K4ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K4ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K4ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K4ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K4ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K4ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K4ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K4ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K4ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K4ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K4ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K4ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K4ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K4ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K4ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K4ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K4ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K4ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K4ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K4ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K4ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K4ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K4ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K4ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K4ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K4ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K4ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K4ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K4ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K4ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K4ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K4ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K4ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K4ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K4ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K4ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K4ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K4ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K4ubuK5}�(K j  )��}�(j�  K j  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K5ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubKj  )��}�(j�  Kj  ]�j�  j�  j  K5ubK j  )��}�(j�  K j  ]�j�  j�  j  K5ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K5ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K5ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K5ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K5ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K5ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K5ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K5ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K5ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K5ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K5ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K5ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K5ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K5ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K5ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K5ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K5ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K5ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K5ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K5ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K5ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K5ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K5ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K5ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K5ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K5ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K5ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K5ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K5ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K5ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K5ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K5ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K5ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K5ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K5ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K5ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K5ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K5ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K5ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K5ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K5ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K5ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K5ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K5ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K5ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K5ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K5ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K5ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K5ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K5ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K5ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K5ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K5ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K5ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K5ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K5ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K5ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K5ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K5ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K5ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K5ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K5ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K5ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K5ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K5ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K5ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K5ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K5ubuK6}�(K j  )��}�(j�  K j  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K6ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubKj  )��}�(j�  Kj  ]�j�  j�  j  K6ubK j  )��}�(j�  K j  ]�j�  j�  j  K6ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K6ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K6ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K6ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K6ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K6ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K6ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K6ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K6ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K6ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K6ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K6ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K6ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K6ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K6ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K6ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K6ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K6ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K6ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K6ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K6ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K6ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K6ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K6ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K6ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K6ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K6ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K6ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K6ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K6ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K6ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K6ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K6ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K6ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K6ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K6ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K6ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K6ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K6ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K6ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K6ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K6ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K6ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K6ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K6ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K6ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K6ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K6ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K6ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K6ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K6ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K6ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K6ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K6ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K6ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K6ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K6ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K6ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K6ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K6ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K6ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K6ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K6ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K6ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K6ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K6ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K6ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K6ubuK7}�(K j  )��}�(j�  K j  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K7ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubKj  )��}�(j�  Kj  ]�j�  j�  j  K7ubK j  )��}�(j�  K j  ]�j�  j�  j  K7ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K7ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K7ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K7ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K7ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K7ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K7ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K7ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K7ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K7ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K7ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K7ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K7ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K7ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K7ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K7ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K7ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K7ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K7ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K7ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K7ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K7ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K7ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K7ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K7ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K7ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K7ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K7ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K7ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K7ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K7ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K7ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K7ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K7ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K7ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K7ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K7ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K7ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K7ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K7ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K7ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K7ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K7ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K7ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K7ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K7ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K7ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K7ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K7ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K7ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K7ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K7ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K7ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K7ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K7ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K7ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K7ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K7ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K7ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K7ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K7ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K7ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K7ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K7ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K7ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K7ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K7ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K7ubuK8}�(K j  )��}�(j�  K j  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K8ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubKj  )��}�(j�  Kj  ]�j�  j�  j  K8ubK j  )��}�(j�  K j  ]�j�  j�  j  K8ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K8ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K8ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K8ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K8ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K8ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K8ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K8ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K8ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K8ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K8ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K8ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K8ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K8ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K8ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K8ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K8ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K8ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K8ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K8ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K8ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K8ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K8ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K8ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K8ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K8ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K8ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K8ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K8ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K8ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K8ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K8ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K8ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K8ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K8ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K8ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K8ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K8ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K8ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K8ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K8ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K8ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K8ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K8ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K8ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K8ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K8ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K8ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K8ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K8ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K8ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K8ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K8ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K8ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K8ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K8ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K8ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K8ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K8ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K8ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K8ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K8ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K8ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K8ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K8ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K8ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K8ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K8ubuK9}�(K j  )��}�(j�  K j  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�K?aj�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�K@aj�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K9ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubKj  )��}�(j�  Kj  ]�j�  j�  j  K9ubK j  )��}�(j�  K j  ]�j�  j�  j  K9ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K9ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K9ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K9ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K9ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K9ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K9ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K9ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K9ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K9ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K9ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K9ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K9ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K9ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K9ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K9ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K9ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K9ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K9ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K9ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K9ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K9ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K9ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K9ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K9ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K9ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K9ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K9ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K9ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K9ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K9ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K9ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K9ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K9ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K9ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K9ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K9ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K9ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K9ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K9ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K9ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K9ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K9ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K9ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K9ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K9ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K9ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K9ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K9ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K9ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K9ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K9ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K9ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K9ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K9ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K9ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K9ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K9ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K9ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K9ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K9ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K9ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K9ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K9ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K9ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K9ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K9ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K9ubuK:}�(K j  )��}�(j�  K j  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K:ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�j�  j�  j  K:ubKj  )��}�(j�  Kj  ]�KCaj�  j�  j  K:ubK j  )��}�(j�  K j  ]�j�  j�  j  K:ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K:ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K:ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K:ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K:ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K:ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K:ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K:ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K:ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K:ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K:ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K:ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K:ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K:ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K:ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K:ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K:ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K:ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K:ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K:ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K:ubK5j  )��}�(j�  K5j  ]��      j�  j�  j  K:ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K:ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K:ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K:ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K:ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K:ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K:ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K:ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K:ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K:ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K:ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K:ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K:ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K:ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K:ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K:ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K:ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K:ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K:ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K:ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K:ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K:ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K:ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K:ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K:ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K:ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K:ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K:ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K:ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K:ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K:ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K:ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K:ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K:ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K:ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K:ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K:ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K:ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K:ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K:ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K:ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K:ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K:ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K:ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K:ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K:ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K:ubuK;}�(K j  )��}�(j�  K j  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K;ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubKj  )��}�(j�  Kj  ]�j�  j�  j  K;ubK j  )��}�(j�  K j  ]�j�  j�  j  K;ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K;ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K;ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K;ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K;ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K;ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K;ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K;ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K;ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K;ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K;ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K;ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K;ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K;ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K;ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K;ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K;ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K;ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K;ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K;ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K;ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K;ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K;ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K;ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K;ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K;ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K;ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K;ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K;ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K;ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K;ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K;ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K;ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K;ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K;ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K;ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K;ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K;ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K;ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K;ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K;ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K;ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K;ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K;ubKLj  )��}�(j�  KLj  ]�KDaj�  j�  j  K;ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K;ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K;ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K;ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K;ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K;ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K;ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K;ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K;ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K;ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K;ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K;ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K;ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K;ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K;ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K;ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K;ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K;ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K;ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K;ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K;ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K;ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K;ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K;ubuK<}�(K j  )��}�(j�  K j  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K<ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubKj  )��}�(j�  Kj  ]�j�  j�  j  K<ubK j  )��}�(j�  K j  ]�j�  j�  j  K<ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K<ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K<ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K<ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K<ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K<ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K<ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K<ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K<ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K<ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K<ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K<ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K<ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K<ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K<ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K<ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K<ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K<ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K<ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K<ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K<ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K<ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K<ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K<ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K<ubK9j  )��}�(j�  K9j  ]�KEaj�  j�  j  K<ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K<ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K<ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K<ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K<ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K<ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K<ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K<ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K<ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K<ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K<ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K<ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K<ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K<ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K<ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K<ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K<ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K<ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K<ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K<ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K<ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K<ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K<ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K<ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K<ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K<ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K<ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K<ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K<ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K<ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K<ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K<ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K<ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K<ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K<ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K<ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K<ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K<ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K<ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K<ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K<ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K<ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K<ubuK=}�(K j  )��}�(j�  K j  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K=ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�j�  j�  j  K=ubKj  )��}�(j�  Kj  ]�KHaj�  j�  j  K=ubK j  )��}�(j�  K j  ]�j�  j�  j  K=ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K=ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K=ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K=ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K=ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K=ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K=ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K=ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K=ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K=ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K=ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K=ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K=ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K=ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K=ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K=ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K=ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K=ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K=ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K=ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K=ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K=ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K=ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K=ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K=ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K=ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K=ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K=ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K=ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K=ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K=ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K=ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K=ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K=ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K=ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K=ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K=ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K=ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K=ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K=ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K=ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K=ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K=ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K=ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K=ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K=ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K=ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K=ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K=ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K=ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K=ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K=ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K=ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K=ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K=ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K=ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K=ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K=ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K=ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K=ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K=ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K=ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K=ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K=ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K=ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K=ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K=ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K=ubuK>}�(K j  )��}�(j�  K j  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�KBaj�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K>ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubKj  )��}�(j�  Kj  ]�j�  j�  j  K>ubK j  )��}�(j�  K j  ]�j�  j�  j  K>ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K>ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K>ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K>ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K>ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K>ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K>ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K>ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K>ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K>ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K>ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K>ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K>ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K>ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K>ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K>ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K>ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K>ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K>ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K>ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K>ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K>ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K>ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K>ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K>ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K>ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K>ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K>ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K>ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K>ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K>ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K>ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K>ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K>ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K>ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K>ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K>ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K>ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K>ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K>ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K>ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K>ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K>ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K>ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K>ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K>ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K>ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K>ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K>ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K>ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K>ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K>ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K>ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K>ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K>ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K>ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K>ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K>ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K>ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K>ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K>ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K>ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K>ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K>ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K>ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K>ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K>ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K>ubuK?}�(K j  )��}�(j�  K j  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�K9aj�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K?ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�j�  j�  j  K?ubKj  )��}�(j�  Kj  ]�KLaj�  j�  j  K?ubK j  )��}�(j�  K j  ]�j�  j�  j  K?ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K?ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K?ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K?ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K?ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K?ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K?ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K?ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K?ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K?ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K?ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K?ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K?ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K?ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K?ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K?ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K?ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K?ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K?ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K?ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K?ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K?ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K?ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K?ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K?ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K?ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K?ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K?ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K?ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K?ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K?ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K?ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K?ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K?ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K?ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K?ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K?ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K?ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K?ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K?ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K?ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K?ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K?ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K?ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K?ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K?ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K?ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K?ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K?ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K?ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K?ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K?ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K?ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K?ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K?ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K?ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K?ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K?ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K?ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K?ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K?ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K?ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K?ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K?ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K?ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K?ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K?ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K?ubuK@}�(K j  )��}�(j�  K j  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K@ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubKj  )��}�(j�  Kj  ]�j�  j�  j  K@ubK j  )��}�(j�  K j  ]�j�  j�  j  K@ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K@ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K@ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K@ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K@ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K@ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K@ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K@ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K@ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K@ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K@ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K@ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K@ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K@ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K@ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K@ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K@ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K@ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K@ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K@ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K@ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K@ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K@ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K@ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K@ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K@ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K@ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K@ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K@ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K@ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K@ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K@ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K@ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K@ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K@ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K@ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K@ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K@ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K@ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K@ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K@ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K@ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K@ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K@ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K@ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K@ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K@ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K@ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K@ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K@ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K@ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K@ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K@ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K@ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K@ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K@ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K@ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K@ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K@ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K@ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K@ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K@ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K@ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K@ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K@ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K@ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K@ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K@ubuKA}�(K j  )��}�(j�  K j  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubK	j  )��}�(j�  K	j  ]�j�  j�  j  KAubK
j  )��}�(j�  K
j  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubKj  )��}�(j�  Kj  ]�j�  j�  j  KAubK j  )��}�(j�  K j  ]�j�  j�  j  KAubK!j  )��}�(j�  K!j  ]�j�  j�  j  KAubK"j  )��}�(j�  K"j  ]�j�  j�  j  KAubK#j  )��}�(j�  K#j  ]�j�  j�  j  KAubK$j  )��}�(j�  K$j  ]�j�  j�  j  KAubK%j  )��}�(j�  K%j  ]�j�  j�  j  KAubK&j  )��}�(j�  K&j  ]�j�  j�  j  KAubK'j  )��}�(j�  K'j  ]�j�  j�  j  KAubK(j  )��}�(j�  K(j  ]�j�  j�  j  KAubK)j  )��}�(j�  K)j  ]�j�  j�  j  KAubK*j  )��}�(j�  K*j  ]�j�  j�  j  KAubK+j  )��}�(j�  K+j  ]�j�  j�  j  KAubK,j  )��}�(j�  K,j  ]�j�  j�  j  KAubK-j  )��}�(j�  K-j  ]�j�  j�  j  KAubK.j  )��}�(j�  K.j  ]�j�  j�  j  KAubK/j  )��}�(j�  K/j  ]�j�  j�  j  KAubK0j  )��}�(j�  K0j  ]�j�  j�  j  KAubK1j  )��}�(j�  K1j  ]�j�  j�  j  KAubK2j  )��}�(j�  K2j  ]�j�  j�  j  KAubK3j  )��}�(j�  K3j  ]�j�  j�  j  KAubK4j  )��}�(j�  K4j  ]�j�  j�  j  KAubK5j  )��}�(j�  K5j  ]�j�  j�  j  KAubK6j  )��}�(j�  K6j  ]�j�  j�  j  KAubK7j  )��}�(j�  K7j  ]�j�  j�  j  KAubK8j  )��}�(j�  K8j  ]�j�  j�  j  KAubK9j  )��}�(j�  K9j  ]�j�  j�  j  KAubK:j  )��}�(j�  K:j  ]�j�  j�  j  KAubK;j  )��}�(j�  K;j  ]�j�  j�  j  KAubK<j  )��}�(j�  K<j  ]�j�  j�  j  KAubK=j  )��}�(j�  K=j  ]�j�  j�  j  KAubK>j  )��}�(j�  K>j  ]�j�  j�  j  KAubK?j  )��}�(j�  K?j  ]�j�  j�  j  KAubK@j  )��}�(j�  K@j  ]�j�  j�  j  KAubKAj  )��}�(j�  KAj  ]�j�  j�  j  KAubKBj  )��}�(j�  KBj  ]�j�  j�  j  KAubKCj  )��}�(j�  KCj  ]�j�  j�  j  KAubKDj  )��}�(j�  KDj  ]�j�  j�  j  KAubKEj  )��}�(j�  KEj  ]�j�  j�  j  KAubKFj  )��}�(j�  KFj  ]�j�  j�  j  KAubKGj  )��}�(j�  KGj  ]�j�  j�  j  KAubKHj  )��}�(j�  KHj  ]�j�  j�  j  KAubKIj  )��}�(j�  KIj  ]�j�  j�  j  KAubKJj  )��}�(j�  KJj  ]�j�  j�  j  KAubKKj  )��}�(j�  KKj  ]�j�  j�  j  KAubKLj  )��}�(j�  KLj  ]�j�  j�  j  KAubKMj  )��}�(j�  KMj  ]�j�  j�  j  KAubKNj  )��}�(j�  KNj  ]�j�  j�  j  KAubKOj  )��}�(j�  KOj  ]�j�  j�  j  KAubKPj  )��}�(j�  KPj  ]�j�  j�  j  KAubKQj  )��}�(j�  KQj  ]�j�  j�  j  KAubKRj  )��}�(j�  KRj  ]�j�  j�  j  KAubKSj  )��}�(j�  KSj  ]�j�  j�  j  KAubKTj  )��}�(j�  KTj  ]�j�  j�  j  KAubKUj  )��}�(j�  KUj  ]�j�  j�  j  KAubKVj  )��}�(j�  KVj  ]�j�  j�  j  KAubKWj  )��}�(j�  KWj  ]�j�  j�  j  KAubKXj  )��}�(j�  KXj  ]�j�  j�  j  KAubKYj  )��}�(j�  KYj  ]�j�  j�  j  KAubKZj  )��}�(j�  KZj  ]�j�  j�  j  KAubK[j  )��}�(j�  K[j  ]�j�  j�  j  KAubK\j  )��}�(j�  K\j  ]�j�  j�  j  KAubK]j  )��}�(j�  K]j  ]�j�  j�  j  KAubK^j  )��}�(j�  K^j  ]�j�  j�  j  KAubK_j  )��}�(j�  K_j  ]�j�  j�  j  KAubK`j  )��}�(j�  K`j  ]�j�  j�  j  KAubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KAubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KAubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KAubuKB}�(K j  )��}�(j�  K j  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�K.aj�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubK	j  )��}�(j�  K	j  ]�j�  j�  j  KBubK
j  )��}�(j�  K
j  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubKj  )��}�(j�  Kj  ]�j�  j�  j  KBubK j  )��}�(j�  K j  ]�j�  j�  j  KBubK!j  )��}�(j�  K!j  ]�j�  j�  j  KBubK"j  )��}�(j�  K"j  ]�j�  j�  j  KBubK#j  )��}�(j�  K#j  ]�j�  j�  j  KBubK$j  )��}�(j�  K$j  ]�j�  j�  j  KBubK%j  )��}�(j�  K%j  ]�j�  j�  j  KBubK&j  )��}�(j�  K&j  ]�j�  j�  j  KBubK'j  )��}�(j�  K'j  ]�j�  j�  j  KBubK(j  )��}�(j�  K(j  ]�j�  j�  j  KBubK)j  )��}�(j�  K)j  ]�j�  j�  j  KBubK*j  )��}�(j�  K*j  ]�j�  j�  j  KBubK+j  )��}�(j�  K+j  ]�j�  j�  j  KBubK,j  )��}�(j�  K,j  ]�j�  j�  j  KBubK-j  )��}�(j�  K-j  ]�j�  j�  j  KBubK.j  )��}�(j�  K.j  ]�j�  j�  j  KBubK/j  )��}�(j�  K/j  ]�j�  j�  j  KBubK0j  )��}�(j�  K0j  ]�j�  j�  j  KBubK1j  )��}�(j�  K1j  ]�j�  j�  j  KBubK2j  )��}�(j�  K2j  ]�j�  j�  j  KBubK3j  )��}�(j�  K3j  ]�j�  j�  j  KBubK4j  )��}�(j�  K4j  ]�j�  j�  j  KBubK5j  )��}�(j�  K5j  ]�j�  j�  j  KBubK6j  )��}�(j�  K6j  ]�j�  j�  j  KBubK7j  )��}�(j�  K7j  ]�j�  j�  j  KBubK8j  )��}�(j�  K8j  ]�j�  j�  j  KBubK9j  )��}�(j�  K9j  ]�j�  j�  j  KBubK:j  )��}�(j�  K:j  ]�j�  j�  j  KBubK;j  )��}�(j�  K;j  ]�j�  j�  j  KBubK<j  )��}�(j�  K<j  ]�j�  j�  j  KBubK=j  )��}�(j�  K=j  ]�j�  j�  j  KBubK>j  )��}�(j�  K>j  ]�j�  j�  j  KBubK?j  )��}�(j�  K?j  ]�j�  j�  j  KBubK@j  )��}�(j�  K@j  ]�j�  j�  j  KBubKAj  )��}�(j�  KAj  ]�j�  j�  j  KBubKBj  )��}�(j�  KBj  ]�j�  j�  j  KBubKCj  )��}�(j�  KCj  ]�j�  j�  j  KBubKDj  )��}�(j�  KDj  ]�j�  j�  j  KBubKEj  )��}�(j�  KEj  ]�j�  j�  j  KBubKFj  )��}�(j�  KFj  ]�j�  j�  j  KBubKGj  )��}�(j�  KGj  ]�j�  j�  j  KBubKHj  )��}�(j�  KHj  ]�j�  j�  j  KBubKIj  )��}�(j�  KIj  ]�j�  j�  j  KBubKJj  )��}�(j�  KJj  ]�j�  j�  j  KBubKKj  )��}�(j�  KKj  ]�j�  j�  j  KBubKLj  )��}�(j�  KLj  ]�j�  j�  j  KBubKMj  )��}�(j�  KMj  ]�j�  j�  j  KBubKNj  )��}�(j�  KNj  ]�j�  j�  j  KBubKOj  )��}�(j�  KOj  ]�j�  j�  j  KBubKPj  )��}�(j�  KPj  ]�j�  j�  j  KBubKQj  )��}�(j�  KQj  ]�j�  j�  j  KBubKRj  )��}�(j�  KRj  ]�j�  j�  j  KBubKSj  )��}�(j�  KSj  ]�j�  j�  j  KBubKTj  )��}�(j�  KTj  ]�j�  j�  j  KBubKUj  )��}�(j�  KUj  ]�j�  j�  j  KBubKVj  )��}�(j�  KVj  ]�j�  j�  j  KBubKWj  )��}�(j�  KWj  ]�j�  j�  j  KBubKXj  )��}�(j�  KXj  ]�j�  j�  j  KBubKYj  )��}�(j�  KYj  ]�j�  j�  j  KBubKZj  )��}�(j�  KZj  ]�j�  j�  j  KBubK[j  )��}�(j�  K[j  ]�j�  j�  j  KBubK\j  )��}�(j�  K\j  ]�j�  j�  j  KBubK]j  )��}�(j�  K]j  ]�j�  j�  j  KBubK^j  )��}�(j�  K^j  ]�j�  j�  j  KBubK_j  )��}�(j�  K_j  ]�j�  j�  j  KBubK`j  )��}�(j�  K`j  ]�j�  j�  j  KBubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KBubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KBubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KBubuKC}�(K j  )��}�(j�  K j  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubK	j  )��}�(j�  K	j  ]�j�  j�  j  KCubK
j  )��}�(j�  K
j  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubKj  )��}�(j�  Kj  ]�j�  j�  j  KCubK j  )��}�(j�  K j  ]�j�  j�  j  KCubK!j  )��}�(j�  K!j  ]�j�  j�  j  KCubK"j  )��}�(j�  K"j  ]�j�  j�  j  KCubK#j  )��}�(j�  K#j  ]�j�  j�  j  KCubK$j  )��}�(j�  K$j  ]�j�  j�  j  KCubK%j  )��}�(j�  K%j  ]�j�  j�  j  KCubK&j  )��}�(j�  K&j  ]�j�  j�  j  KCubK'j  )��}�(j�  K'j  ]�j�  j�  j  KCubK(j  )��}�(j�  K(j  ]�j�  j�  j  KCubK)j  )��}�(j�  K)j  ]�j�  j�  j  KCubK*j  )��}�(j�  K*j  ]�j�  j�  j  KCubK+j  )��}�(j�  K+j  ]�j�  j�  j  KCubK,j  )��}�(j�  K,j  ]�j�  j�  j  KCubK-j  )��}�(j�  K-j  ]�j�  j�  j  KCubK.j  )��}�(j�  K.j  ]�j�  j�  j  KCubK/j  )��}�(j�  K/j  ]�j�  j�  j  KCubK0j  )��}�(j�  K0j  ]�j�  j�  j  KCubK1j  )��}�(j�  K1j  ]�j�  j�  j  KCubK2j  )��}�(j�  K2j  ]�j�  j�  j  KCubK3j  )��}�(j�  K3j  ]�j�  j�  j  KCubK4j  )��}�(j�  K4j  ]�j�  j�  j  KCubK5j  )��}�(j�  K5j  ]�j�  j�  j  KCubK6j  )��}�(j�  K6j  ]�j�  j�  j  KCubK7j  )��}�(j�  K7j  ]�j�  j�  j  KCubK8j  )��}�(j�  K8j  ]�j�  j�  j  KCubK9j  )��}�(j�  K9j  ]�j�  j�  j  KCubK:j  )��}�(j�  K:j  ]�j�  j�  j  KCubK;j  )��}�(j�  K;j  ]�j�  j�  j  KCubK<j  )��}�(j�  K<j  ]�j�  j�  j  KCubK=j  )��}�(j�  K=j  ]�j�  j�  j  KCubK>j  )��}�(j�  K>j  ]�j�  j�  j  KCubK?j  )��}�(j�  K?j  ]�j�  j�  j  KCubK@j  )��}�(j�  K@j  ]�j�  j�  j  KCubKAj  )��}�(j�  KAj  ]�j�  j�  j  KCubKBj  )��}�(j�  KBj  ]�j�  j�  j  KCubKCj  )��}�(j�  KCj  ]�j�  j�  j  KCubKDj  )��}�(j�  KDj  ]�j�  j�  j  KCubKEj  )��}�(j�  KEj  ]�j�  j�  j  KCubKFj  )��}�(j�  KFj  ]�j�  j�  j  KCubKGj  )��}�(j�  KGj  ]�j�  j�  j  KCubKHj  )��}�(j�  KHj  ]�j�  j�  j  KCubKIj  )��}�(j�  KIj  ]�j�  j�  j  KCubKJj  )��}�(j�  KJj  ]�j�  j�  j  KCubKKj  )��}�(j�  KKj  ]�j�  j�  j  KCubKLj  )��}�(j�  KLj  ]�j�  j�  j  KCubKMj  )��}�(j�  KMj  ]�j�  j�  j  KCubKNj  )��}�(j�  KNj  ]�j�  j�  j  KCubKOj  )��}�(j�  KOj  ]�j�  j�  j  KCubKPj  )��}�(j�  KPj  ]�j�  j�  j  KCubKQj  )��}�(j�  KQj  ]�j�  j�  j  KCubKRj  )��}�(j�  KRj  ]�j�  j�  j  KCubKSj  )��}�(j�  KSj  ]�j�  j�  j  KCubKTj  )��}�(j�  KTj  ]�j�  j�  j  KCubKUj  )��}�(j�  KUj  ]�j�  j�  j  KCubKVj  )��}�(j�  KVj  ]�j�  j�  j  KCubKWj  )��}�(j�  KWj  ]�j�  j�  j  KCubKXj  )��}�(j�  KXj  ]�j�  j�  j  KCubKYj  )��}�(j�  KYj  ]�j�  j�  j  KCubKZj  )��}�(j�  KZj  ]�j�  j�  j  KCubK[j  )��}�(j�  K[j  ]�j�  j�  j  KCubK\j  )��}�(j�  K\j  ]�j�  j�  j  KCubK]j  )��}�(j�  K]j  ]�j�  j�  j  KCubK^j  )��}�(j�  K^j  ]�j�  j�  j  KCubK_j  )��}�(j�  K_j  ]�j�  j�  j  KCubK`j  )��}�(j�  K`j  ]�j�  j�  j  KCubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KCubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KCubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KCubuKD}�(K j  )��}�(j�  K j  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubK	j  )��}�(j�  K	j  ]�j�  j�  j  KDubK
j  )��}�(j�  K
j  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubKj  )��}�(j�  Kj  ]�j�  j�  j  KDubK j  )��}�(j�  K j  ]�j�  j�  j  KDubK!j  )��}�(j�  K!j  ]�j�  j�  j  KDubK"j  )��}�(j�  K"j  ]�j�  j�  j  KDubK#j  )��}�(j�  K#j  ]�j�  j�  j  KDubK$j  )��}�(j�  K$j  ]�j�  j�  j  KDubK%j  )��}�(j�  K%j  ]�j�  j�  j  KDubK&j  )��}�(j�  K&j  ]�j�  j�  j  KDubK'j  )��}�(j�  K'j  ]�j�  j�  j  KDubK(j  )��}�(j�  K(j  ]�j�  j�  j  KDubK)j  )��}�(j�  K)j  ]�j�  j�  j  KDubK*j  )��}�(j�  K*j  ]�j�  j�  j  KDubK+j  )��}�(j�  K+j  ]�j�  j�  j  KDubK,j  )��}�(j�  K,j  ]�j�  j�  j  KDubK-j  )��}�(j�  K-j  ]�j�  j�  j  KDubK.j  )��}�(j�  K.j  ]�j�  j�  j  KDubK/j  )��}�(j�  K/j  ]�j�  j�  j  KDubK0j  )��}�(j�  K0j  ]�j�  j�  j  KDubK1j  )��}�(j�  K1j  ]�j�  j�  j  KDubK2j  )��}�(j�  K2j  ]�j�  j�  j  KDubK3j  )��}�(j�  K3j  ]�j�  j�  j  KDubK4j  )��}�(j�  K4j  ]�j�  j�  j  KDubK5j  )��}�(j�  K5j  ]�j�  j�  j  KDubK6j  )��}�(j�  K6j  ]�j�  j�  j  KDubK7j  )��}�(j�  K7j  ]�j�  j�  j  KDubK8j  )��}�(j�  K8j  ]�j�  j�  j  KDubK9j  )��}�(j�  K9j  ]�j�  j�  j  KDubK:j  )��}�(j�  K:j  ]�j�  j�  j  KDubK;j  )��}�(j�  K;j  ]�j�  j�  j  KDubK<j  )��}�(j�  K<j  ]�j�  j�  j  KDubK=j  )��}�(j�  K=j  ]�j�  j�  j  KDubK>j  )��}�(j�  K>j  ]�j�  j�  j  KDubK?j  )��}�(j�  K?j  ]�j�  j�  j  KDubK@j  )��}�(j�  K@j  ]�j�  j�  j  KDubKAj  )��}�(j�  KAj  ]�j�  j�  j  KDubKBj  )��}�(j�  KBj  ]�j�  j�  j  KDubKCj  )��}�(j�  KCj  ]�j�  j�  j  KDubKDj  )��}�(j�  KDj  ]�j�  j�  j  KDubKEj  )��}�(j�  KEj  ]�j�  j�  j  KDubKFj  )��}�(j�  KFj  ]�j�  j�  j  KDubKGj  )��}�(j�  KGj  ]�j�  j�  j  KDubKHj  )��}�(j�  KHj  ]�j�  j�  j  KDubKIj  )��}�(j�  KIj  ]�j�  j�  j  KDubKJj  )��}�(j�  KJj  ]�j�  j�  j  KDubKKj  )��}�(j�  KKj  ]�j�  j�  j  KDubKLj  )��}�(j�  KLj  ]�j�  j�  j  KDubKMj  )��}�(j�  KMj  ]�j�  j�  j  KDubKNj  )��}�(j�  KNj  ]�j�  j�  j  KDubKOj  )��}�(j�  KOj  ]�j�  j�  j  KDubKPj  )��}�(j�  KPj  ]�j�  j�  j  KDubKQj  )��}�(j�  KQj  ]�j�  j�  j  KDubKRj  )��}�(j�  KRj  ]�j�  j�  j  KDubKSj  )��}�(j�  KSj  ]�j�  j�  j  KDubKTj  )��}�(j�  KTj  ]�j�  j�  j  KDubKUj  )��}�(j�  KUj  ]�j�  j�  j  KDubKVj  )��}�(j�  KVj  ]�j�  j�  j  KDubKWj  )��}�(j�  KWj  ]�j�  j�  j  KDubKXj  )��}�(j�  KXj  ]�j�  j�  j  KDubKYj  )��}�(j�  KYj  ]�j�  j�  j  KDubKZj  )��}�(j�  KZj  ]�j�  j�  j  KDubK[j  )��}�(j�  K[j  ]�j�  j�  j  KDubK\j  )��}�(j�  K\j  ]�j�  j�  j  KDubK]j  )��}�(j�  K]j  ]�j�  j�  j  KDubK^j  )��}�(j�  K^j  ]�j�  j�  j  KDubK_j  )��}�(j�  K_j  ]�j�  j�  j  KDubK`j  )��}�(j�  K`j  ]�j�  j�  j  KDubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KDubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KDubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KDubuKE}�(K j  )��}�(j�  K j  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�KKaj�  j�  j  KEubKj  )��}�(j�  Kj  ]�KWaj�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�KPaj�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubK	j  )��}�(j�  K	j  ]�j�  j�  j  KEubK
j  )��}�(j�  K
j  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubKj  )��}�(j�  Kj  ]�j�  j�  j  KEubK j  )��}�(j�  K j  ]�j�  j�  j  KEubK!j  )��}�(j�  K!j  ]�j�  j�  j  KEubK"j  )��}�(j�  K"j  ]�j�  j�  j  KEubK#j  )��}�(j�  K#j  ]�j�  j�  j  KEubK$j  )��}�(j�  K$j  ]�j�  j�  j  KEubK%j  )��}�(j�  K%j  ]�j�  j�  j  KEubK&j  )��}�(j�  K&j  ]�j�  j�  j  KEubK'j  )��}�(j�  K'j  ]�j�  j�  j  KEubK(j  )��}�(j�  K(j  ]�j�  j�  j  KEubK)j  )��}�(j�  K)j  ]�j�  j�  j  KEubK*j  )��}�(j�  K*j  ]�j�  j�  j  KEubK+j  )��}�(j�  K+j  ]�j�  j�  j  KEubK,j  )��}�(j�  K,j  ]�j�  j�  j  KEubK-j  )��}�(j�  K-j  ]�j�  j�  j  KEubK.j  )��}�(j�  K.j  ]�j�  j�  j  KEubK/j  )��}�(j�  K/j  ]�j�  j�  j  KEubK0j  )��}�(j�  K0j  ]�j�  j�  j  KEubK1j  )��}�(j�  K1j  ]�j�  j�  j  KEubK2j  )��}�(j�  K2j  ]�j�  j�  j  KEubK3j  )��}�(j�  K3j  ]�j�  j�  j  KEubK4j  )��}�(j�  K4j  ]�j�  j�  j  KEubK5j  )��}�(j�  K5j  ]�j�  j�  j  KEubK6j  )��}�(j�  K6j  ]�j�  j�  j  KEubK7j  )��}�(j�  K7j  ]�j�  j�  j  KEubK8j  )��}�(j�  K8j  ]�j�  j�  j  KEubK9j  )��}�(j�  K9j  ]�j�  j�  j  KEubK:j  )��}�(j�  K:j  ]�j�  j�  j  KEubK;j  )��}�(j�  K;j  ]�j�  j�  j  KEubK<j  )��}�(j�  K<j  ]�j�  j�  j  KEubK=j  )��}�(j�  K=j  ]�j�  j�  j  KEubK>j  )��}�(j�  K>j  ]�j�  j�  j  KEubK?j  )��}�(j�  K?j  ]�j�  j�  j  KEubK@j  )��}�(j�  K@j  ]�j�  j�  j  KEubKAj  )��}�(j�  KAj  ]�j�  j�  j  KEubKBj  )��}�(j�  KBj  ]�j�  j�  j  KEubKCj  )��}�(j�  KCj  ]�j�  j�  j  KEubKDj  )��}�(j�  KDj  ]�j�  j�  j  KEubKEj  )��}�(j�  KEj  ]�j�  j�  j  KEubKFj  )��}�(j�  KFj  ]�j�  j�  j  KEubKGj  )��}�(j�  KGj  ]�j�  j�  j  KEubKHj  )��}�(j�  KHj  ]�j�  j�  j  KEubKIj  )��}�(j�  KIj  ]�j�  j�  j  KEubKJj  )��}�(j�  KJj  ]�j�  j�  j  KEubKKj  )��}�(j�  KKj  ]�j�  j�  j  KEubKLj  )��}�(j�  KLj  ]�j�  j�  j  KEubKMj  )��}�(j�  KMj  ]�j�  j�  j  KEubKNj  )��}�(j�  KNj  ]�j�  j�  j  KEubKOj  )��}�(j�  KOj  ]�j�  j�  j  KEubKPj  )��}�(j�  KPj  ]�j�  j�  j  KEubKQj  )��}�(j�  KQj  ]�j�  j�  j  KEubKRj  )��}�(j�  KRj  ]�j�  j�  j  KEubKSj  )��}�(j�  KSj  ]�j�  j�  j  KEubKTj  )��}�(j�  KTj  ]�j�  j�  j  KEubKUj  )��}�(j�  KUj  ]�j�  j�  j  KEubKVj  )��}�(j�  KVj  ]�j�  j�  j  KEubKWj  )��}�(j�  KWj  ]�j�  j�  j  KEubKXj  )��}�(j�  KXj  ]�j�  j�  j  KEubKYj  )��}�(j�  KYj  ]�j�  j�  j  KEubKZj  )��}�(j�  KZj  ]�j�  j�  j  KEubK[j  )��}�(j�  K[j  ]�j�  j�  j  KEubK\j  )��}�(j�  K\j  ]�j�  j�  j  KEubK]j  )��}�(j�  K]j  ]�j�  j�  j  KEubK^j  )��}�(j�  K^j  ]�j�  j�  j  KEubK_j  )��}�(j�  K_j  ]�j�  j�  j  KEubK`j  )��}�(j�  K`j  ]�j�  j�  j  KEubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KEubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KEubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KEubuKF}�(K j  )��}�(j�  K j  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubK	j  )��}�(j�  K	j  ]�j�  j�  j  KFubK
j  )��}�(j�  K
j  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubKj  )��}�(j�  Kj  ]�j�  j�  j  KFubK j  )��}�(j�  K j  ]�j�  j�  j  KFubK!j  )��}�(j�  K!j  ]�j�  j�  j  KFubK"j  )��}�(j�  K"j  ]�j�  j�  j  KFubK#j  )��}�(j�  K#j  ]�j�  j�  j  KFubK$j  )��}�(j�  K$j  ]�j�  j�  j  KFubK%j  )��}�(j�  K%j  ]�j�  j�  j  KFubK&j  )��}�(j�  K&j  ]�j�  j�  j  KFubK'j  )��}�(j�  K'j  ]�j�  j�  j  KFubK(j  )��}�(j�  K(j  ]�j�  j�  j  KFubK)j  )��}�(j�  K)j  ]�j�  j�  j  KFubK*j  )��}�(j�  K*j  ]�j�  j�  j  KFubK+j  )��}�(j�  K+j  ]�j�  j�  j  KFubK,j  )��}�(j�  K,j  ]�j�  j�  j  KFubK-j  )��}�(j�  K-j  ]�j�  j�  j  KFubK.j  )��}�(j�  K.j  ]�j�  j�  j  KFubK/j  )��}�(j�  K/j  ]�j�  j�  j  KFubK0j  )��}�(j�  K0j  ]�j�  j�  j  KFubK1j  )��}�(j�  K1j  ]�j�  j�  j  KFubK2j  )��}�(j�  K2j  ]�j�  j�  j  KFubK3j  )��}�(j�  K3j  ]�j�  j�  j  KFubK4j  )��}�(j�  K4j  ]�j�  j�  j  KFubK5j  )��}�(j�  K5j  ]�j�  j�  j  KFubK6j  )��}�(j�  K6j  ]�j�  j�  j  KFubK7j  )��}�(j�  K7j  ]�j�  j�  j  KFubK8j  )��}�(j�  K8j  ]�j�  j�  j  KFubK9j  )��}�(j�  K9j  ]�j�  j�  j  KFubK:j  )��}�(j�  K:j  ]�j�  j�  j  KFubK;j  )��}�(j�  K;j  ]�j�  j�  j  KFubK<j  )��}�(j�  K<j  ]�j�  j�  j  KFubK=j  )��}�(j�  K=j  ]�j�  j�  j  KFubK>j  )��}�(j�  K>j  ]�j�  j�  j  KFubK?j  )��}�(j�  K?j  ]�j�  j�  j  KFubK@j  )��}�(j�  K@j  ]�j�  j�  j  KFubKAj  )��}�(j�  KAj  ]�j�  j�  j  KFubKBj  )��}�(j�  KBj  ]�j�  j�  j  KFubKCj  )��}�(j�  KCj  ]�j�  j�  j  KFubKDj  )��}�(j�  KDj  ]�j�  j�  j  KFubKEj  )��}�(j�  KEj  ]�j�  j�  j  KFubKFj  )��}�(j�  KFj  ]�j�  j�  j  KFubKGj  )��}�(j�  KGj  ]�j�  j�  j  KFubKHj  )��}�(j�  KHj  ]�j�  j�  j  KFubKIj  )��}�(j�  KIj  ]�j�  j�  j  KFubKJj  )��}�(j�  KJj  ]�j�  j�  j  KFubKKj  )��}�(j�  KKj  ]�j�  j�  j  KFubKLj  )��}�(j�  KLj  ]�j�  j�  j  KFubKMj  )��}�(j�  KMj  ]�j�  j�  j  KFubKNj  )��}�(j�  KNj  ]�j�  j�  j  KFubKOj  )��}�(j�  KOj  ]�j�  j�  j  KFubKPj  )��}�(j�  KPj  ]�j�  j�  j  KFubKQj  )��}�(j�  KQj  ]�j�  j�  j  KFubKRj  )��}�(j�  KRj  ]�j�  j�  j  KFubKSj  )��}�(j�  KSj  ]�j�  j�  j  KFubKTj  )��}�(j�  KTj  ]�j�  j�  j  KFubKUj  )��}�(j�  KUj  ]�j�  j�  j  KFubKVj  )��}�(j�  KVj  ]�j�  j�  j  KFubKWj  )��}�(j�  KWj  ]�j�  j�  j  KFubKXj  )��}�(j�  KXj  ]�j�  j�  j  KFubKYj  )��}�(j�  KYj  ]�j�  j�  j  KFubKZj  )��}�(j�  KZj  ]�j�  j�  j  KFubK[j  )��}�(j�  K[j  ]�j�  j�  j  KFubK\j  )��}�(j�  K\j  ]�j�  j�  j  KFubK]j  )��}�(j�  K]j  ]�j�  j�  j  KFubK^j  )��}�(j�  K^j  ]�j�  j�  j  KFubK_j  )��}�(j�  K_j  ]�j�  j�  j  KFubK`j  )��}�(j�  K`j  ]�j�  j�  j  KFubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KFubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KFubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KFubuKG}�(K j  )��}�(j�  K j  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�K[aj�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubK	j  )��}�(j�  K	j  ]�j�  j�  j  KGubK
j  )��}�(j�  K
j  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubKj  )��}�(j�  Kj  ]�j�  j�  j  KGubK j  )��}�(j�  K j  ]�j�  j�  j  KGubK!j  )��}�(j�  K!j  ]�j�  j�  j  KGubK"j  )��}�(j�  K"j  ]�j�  j�  j  KGubK#j  )��}�(j�  K#j  ]�j�  j�  j  KGubK$j  )��}�(j�  K$j  ]�j�  j�  j  KGubK%j  )��}�(j�  K%j  ]�j�  j�  j  KGubK&j  )��}�(j�  K&j  ]�j�  j�  j  KGubK'j  )��}�(j�  K'j  ]�j�  j�  j  KGubK(j  )��}�(j�  K(j  ]�j�  j�  j  KGubK)j  )��}�(j�  K)j  ]�j�  j�  j  KGubK*j  )��}�(j�  K*j  ]�j�  j�  j  KGubK+j  )��}�(j�  K+j  ]�j�  j�  j  KGubK,j  )��}�(j�  K,j  ]�j�  j�  j  KGubK-j  )��}�(j�  K-j  ]�j�  j�  j  KGubK.j  )��}�(j�  K.j  ]�j�  j�  j  KGubK/j  )��}�(j�  K/j  ]�j�  j�  j  KGubK0j  )��}�(j�  K0j  ]�j�  j�  j  KGubK1j  )��}�(j�  K1j  ]�j�  j�  j  KGubK2j  )��}�(j�  K2j  ]�j�  j�  j  KGubK3j  )��}�(j�  K3j  ]�j�  j�  j  KGubK4j  )��}�(j�  K4j  ]�j�  j�  j  KGubK5j  )��}�(j�  K5j  ]�j�  j�  j  KGubK6j  )��}�(j�  K6j  ]�j�  j�  j  KGubK7j  )��}�(j�  K7j  ]�j�  j�  j  KGubK8j  )��}�(j�  K8j  ]�j�  j�  j  KGubK9j  )��}�(j�  K9j  ]�j�  j�  j  KGubK:j  )��}�(j�  K:j  ]�j�  j�  j  KGubK;j  )��}�(j�  K;j  ]�j�  j�  j  KGubK<j  )��}�(j�  K<j  ]�j�  j�  j  KGubK=j  )��}�(j�  K=j  ]�j�  j�  j  KGubK>j  )��}�(j�  K>j  ]�j�  j�  j  KGubK?j  )��}�(j�  K?j  ]�j�  j�  j  KGubK@j  )��}�(j�  K@j  ]�j�  j�  j  KGubKAj  )��}�(j�  KAj  ]�j�  j�  j  KGubKBj  )��}�(j�  KBj  ]�j�  j�  j  KGubKCj  )��}�(j�  KCj  ]�j�  j�  j  KGubKDj  )��}�(j�  KDj  ]�j�  j�  j  KGubKEj  )��}�(j�  KEj  ]�j�  j�  j  KGubKFj  )��}�(j�  KFj  ]�j�  j�  j  KGubKGj  )��}�(j�  KGj  ]�j�  j�  j  KGubKHj  )��}�(j�  KHj  ]�j�  j�  j  KGubKIj  )��}�(j�  KIj  ]�j�  j�  j  KGubKJj  )��}�(j�  KJj  ]�j�  j�  j  KGubKKj  )��}�(j�  KKj  ]�j�  j�  j  KGubKLj  )��}�(j�  KLj  ]�j�  j�  j  KGubKMj  )��}�(j�  KMj  ]�j�  j�  j  KGubKNj  )��}�(j�  KNj  ]�j�  j�  j  KGubKOj  )��}�(j�  KOj  ]�j�  j�  j  KGubKPj  )��}�(j�  KPj  ]�j�  j�  j  KGubKQj  )��}�(j�  KQj  ]�j�  j�  j  KGubKRj  )��}�(j�  KRj  ]�j�  j�  j  KGubKSj  )��}�(j�  KSj  ]�j�  j�  j  KGubKTj  )��}�(j�  KTj  ]�j�  j�  j  KGubKUj  )��}�(j�  KUj  ]�j�  j�  j  KGubKVj  )��}�(j�  KVj  ]�j�  j�  j  KGubKWj  )��}�(j�  KWj  ]�j�  j�  j  KGubKXj  )��}�(j�  KXj  ]�j�  j�  j  KGubKYj  )��}�(j�  KYj  ]�j�  j�  j  KGubKZj  )��}�(j�  KZj  ]�j�  j�  j  KGubK[j  )��}�(j�  K[j  ]�j�  j�  j  KGubK\j  )��}�(j�  K\j  ]�j�  j�  j  KGubK]j  )��}�(j�  K]j  ]�j�  j�  j  KGubK^j  )��}�(j�  K^j  ]�j�  j�  j  KGubK_j  )��}�(j�  K_j  ]�j�  j�  j  KGubK`j  )��}�(j�  K`j  ]�j�  j�  j  KGubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KGubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KGubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KGubuKH}�(K j  )��}�(j�  K j  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubK	j  )��}�(j�  K	j  ]�j�  j�  j  KHubK
j  )��}�(j�  K
j  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubKj  )��}�(j�  Kj  ]�j�  j�  j  KHubK j  )��}�(j�  K j  ]�j�  j�  j  KHubK!j  )��}�(j�  K!j  ]�j�  j�  j  KHubK"j  )��}�(j�  K"j  ]�j�  j�  j  KHubK#j  )��}�(j�  K#j  ]�j�  j�  j  KHubK$j  )��}�(j�  K$j  ]�j�  j�  j  KHubK%j  )��}�(j�  K%j  ]�j�  j�  j  KHubK&j  )��}�(j�  K&j  ]�j�  j�  j  KHubK'j  )��}�(j�  K'j  ]�j�  j�  j  KHubK(j  )��}�(j�  K(j  ]�j�  j�  j  KHubK)j  )��}�(j�  K)j  ]�j�  j�  j  KHubK*j  )��}�(j�  K*j  ]�j�  j�  j  KHubK+j  )��}�(j�  K+j  ]�j�  j�  j  KHubK,j  )��}�(j�  K,j  ]�j�  j�  j  KHubK-j  )��}�(j�  K-j  ]�j�  j�  j  KHubK.j  )��}�(j�  K.j  ]�j�  j�  j  KHubK/j  )��}�(j�  K/j  ]�j�  j�  j  KHubK0j  )��}�(j�  K0j  ]�j�  j�  j  KHubK1j  )��}�(j�  K1j  ]�j�  j�  j  KHubK2j  )��}�(j�  K2j  ]�j�  j�  j  KHubK3j  )��}�(j�  K3j  ]�j�  j�  j  KHubK4j  )��}�(j�  K4j  ]�j�  j�  j  KHubK5j  )��}�(j�  K5j  ]�j�  j�  j  KHubK6j  )��}�(j�  K6j  ]�j�  j�  j  KHubK7j  )��}�(j�  K7j  ]�j�  j�  j  KHubK8j  )��}�(j�  K8j  ]�j�  j�  j  KHubK9j  )��}�(j�  K9j  ]�j�  j�  j  KHubK:j  )��}�(j�  K:j  ]�j�  j�  j  KHubK;j  )��}�(j�  K;j  ]�j�  j�  j  KHubK<j  )��}�(j�  K<j  ]�j�  j�  j  KHubK=j  )��}�(j�  K=j  ]�j�  j�  j  KHubK>j  )��}�(j�  K>j  ]�j�  j�  j  KHubK?j  )��}�(j�  K?j  ]�j�  j�  j  KHubK@j  )��}�(j�  K@j  ]�j�  j�  j  KHubKAj  )��}�(j�  KAj  ]�j�  j�  j  KHubKBj  )��}�(j�  KBj  ]�j�  j�  j  KHubKCj  )��}�(j�  KCj  ]�j�  j�  j  KHubKDj  )��}�(j�  KDj  ]�j�  j�  j  KHubKEj  )��}�(j�  KEj  ]�j�  j�  j  KHubKFj  )��}�(j�  KFj  ]�j�  j�  j  KHubKGj  )��}�(j�  KGj  ]�j�  j�  j  KHubKHj  )��}�(j�  KHj  ]�j�  j�  j  KHubKIj  )��}�(j�  KIj  ]�j�  j�  j  KHubKJj  )��}�(j�  KJj  ]�j�  j�  j  KHubKKj  )��}�(j�  KKj  ]�j�  j�  �      j  KHubKLj  )��}�(j�  KLj  ]�j�  j�  j  KHubKMj  )��}�(j�  KMj  ]�j�  j�  j  KHubKNj  )��}�(j�  KNj  ]�j�  j�  j  KHubKOj  )��}�(j�  KOj  ]�j�  j�  j  KHubKPj  )��}�(j�  KPj  ]�j�  j�  j  KHubKQj  )��}�(j�  KQj  ]�j�  j�  j  KHubKRj  )��}�(j�  KRj  ]�j�  j�  j  KHubKSj  )��}�(j�  KSj  ]�j�  j�  j  KHubKTj  )��}�(j�  KTj  ]�j�  j�  j  KHubKUj  )��}�(j�  KUj  ]�j�  j�  j  KHubKVj  )��}�(j�  KVj  ]�j�  j�  j  KHubKWj  )��}�(j�  KWj  ]�j�  j�  j  KHubKXj  )��}�(j�  KXj  ]�j�  j�  j  KHubKYj  )��}�(j�  KYj  ]�j�  j�  j  KHubKZj  )��}�(j�  KZj  ]�j�  j�  j  KHubK[j  )��}�(j�  K[j  ]�j�  j�  j  KHubK\j  )��}�(j�  K\j  ]�j�  j�  j  KHubK]j  )��}�(j�  K]j  ]�j�  j�  j  KHubK^j  )��}�(j�  K^j  ]�j�  j�  j  KHubK_j  )��}�(j�  K_j  ]�j�  j�  j  KHubK`j  )��}�(j�  K`j  ]�j�  j�  j  KHubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KHubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KHubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KHubuKI}�(K j  )��}�(j�  K j  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubK	j  )��}�(j�  K	j  ]�j�  j�  j  KIubK
j  )��}�(j�  K
j  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubKj  )��}�(j�  Kj  ]�j�  j�  j  KIubK j  )��}�(j�  K j  ]�j�  j�  j  KIubK!j  )��}�(j�  K!j  ]�j�  j�  j  KIubK"j  )��}�(j�  K"j  ]�j�  j�  j  KIubK#j  )��}�(j�  K#j  ]�j�  j�  j  KIubK$j  )��}�(j�  K$j  ]�j�  j�  j  KIubK%j  )��}�(j�  K%j  ]�j�  j�  j  KIubK&j  )��}�(j�  K&j  ]�j�  j�  j  KIubK'j  )��}�(j�  K'j  ]�j�  j�  j  KIubK(j  )��}�(j�  K(j  ]�j�  j�  j  KIubK)j  )��}�(j�  K)j  ]�j�  j�  j  KIubK*j  )��}�(j�  K*j  ]�j�  j�  j  KIubK+j  )��}�(j�  K+j  ]�j�  j�  j  KIubK,j  )��}�(j�  K,j  ]�j�  j�  j  KIubK-j  )��}�(j�  K-j  ]�j�  j�  j  KIubK.j  )��}�(j�  K.j  ]�j�  j�  j  KIubK/j  )��}�(j�  K/j  ]�j�  j�  j  KIubK0j  )��}�(j�  K0j  ]�j�  j�  j  KIubK1j  )��}�(j�  K1j  ]�j�  j�  j  KIubK2j  )��}�(j�  K2j  ]�j�  j�  j  KIubK3j  )��}�(j�  K3j  ]�j�  j�  j  KIubK4j  )��}�(j�  K4j  ]�j�  j�  j  KIubK5j  )��}�(j�  K5j  ]�j�  j�  j  KIubK6j  )��}�(j�  K6j  ]�j�  j�  j  KIubK7j  )��}�(j�  K7j  ]�j�  j�  j  KIubK8j  )��}�(j�  K8j  ]�j�  j�  j  KIubK9j  )��}�(j�  K9j  ]�j�  j�  j  KIubK:j  )��}�(j�  K:j  ]�j�  j�  j  KIubK;j  )��}�(j�  K;j  ]�j�  j�  j  KIubK<j  )��}�(j�  K<j  ]�j�  j�  j  KIubK=j  )��}�(j�  K=j  ]�j�  j�  j  KIubK>j  )��}�(j�  K>j  ]�j�  j�  j  KIubK?j  )��}�(j�  K?j  ]�j�  j�  j  KIubK@j  )��}�(j�  K@j  ]�j�  j�  j  KIubKAj  )��}�(j�  KAj  ]�j�  j�  j  KIubKBj  )��}�(j�  KBj  ]�j�  j�  j  KIubKCj  )��}�(j�  KCj  ]�j�  j�  j  KIubKDj  )��}�(j�  KDj  ]�j�  j�  j  KIubKEj  )��}�(j�  KEj  ]�j�  j�  j  KIubKFj  )��}�(j�  KFj  ]�j�  j�  j  KIubKGj  )��}�(j�  KGj  ]�j�  j�  j  KIubKHj  )��}�(j�  KHj  ]�j�  j�  j  KIubKIj  )��}�(j�  KIj  ]�j�  j�  j  KIubKJj  )��}�(j�  KJj  ]�j�  j�  j  KIubKKj  )��}�(j�  KKj  ]�j�  j�  j  KIubKLj  )��}�(j�  KLj  ]�j�  j�  j  KIubKMj  )��}�(j�  KMj  ]�j�  j�  j  KIubKNj  )��}�(j�  KNj  ]�j�  j�  j  KIubKOj  )��}�(j�  KOj  ]�j�  j�  j  KIubKPj  )��}�(j�  KPj  ]�j�  j�  j  KIubKQj  )��}�(j�  KQj  ]�j�  j�  j  KIubKRj  )��}�(j�  KRj  ]�j�  j�  j  KIubKSj  )��}�(j�  KSj  ]�j�  j�  j  KIubKTj  )��}�(j�  KTj  ]�j�  j�  j  KIubKUj  )��}�(j�  KUj  ]�j�  j�  j  KIubKVj  )��}�(j�  KVj  ]�j�  j�  j  KIubKWj  )��}�(j�  KWj  ]�j�  j�  j  KIubKXj  )��}�(j�  KXj  ]�j�  j�  j  KIubKYj  )��}�(j�  KYj  ]�j�  j�  j  KIubKZj  )��}�(j�  KZj  ]�j�  j�  j  KIubK[j  )��}�(j�  K[j  ]�j�  j�  j  KIubK\j  )��}�(j�  K\j  ]�j�  j�  j  KIubK]j  )��}�(j�  K]j  ]�j�  j�  j  KIubK^j  )��}�(j�  K^j  ]�j�  j�  j  KIubK_j  )��}�(j�  K_j  ]�j�  j�  j  KIubK`j  )��}�(j�  K`j  ]�j�  j�  j  KIubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KIubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KIubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KIubuKJ}�(K j  )��}�(j�  K j  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubK	j  )��}�(j�  K	j  ]�j�  j�  j  KJubK
j  )��}�(j�  K
j  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�KMaj�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubKj  )��}�(j�  Kj  ]�j�  j�  j  KJubK j  )��}�(j�  K j  ]�j�  j�  j  KJubK!j  )��}�(j�  K!j  ]�j�  j�  j  KJubK"j  )��}�(j�  K"j  ]�j�  j�  j  KJubK#j  )��}�(j�  K#j  ]�j�  j�  j  KJubK$j  )��}�(j�  K$j  ]�j�  j�  j  KJubK%j  )��}�(j�  K%j  ]�j�  j�  j  KJubK&j  )��}�(j�  K&j  ]�j�  j�  j  KJubK'j  )��}�(j�  K'j  ]�j�  j�  j  KJubK(j  )��}�(j�  K(j  ]�j�  j�  j  KJubK)j  )��}�(j�  K)j  ]�j�  j�  j  KJubK*j  )��}�(j�  K*j  ]�j�  j�  j  KJubK+j  )��}�(j�  K+j  ]�j�  j�  j  KJubK,j  )��}�(j�  K,j  ]�j�  j�  j  KJubK-j  )��}�(j�  K-j  ]�j�  j�  j  KJubK.j  )��}�(j�  K.j  ]�j�  j�  j  KJubK/j  )��}�(j�  K/j  ]�j�  j�  j  KJubK0j  )��}�(j�  K0j  ]�j�  j�  j  KJubK1j  )��}�(j�  K1j  ]�j�  j�  j  KJubK2j  )��}�(j�  K2j  ]�j�  j�  j  KJubK3j  )��}�(j�  K3j  ]�j�  j�  j  KJubK4j  )��}�(j�  K4j  ]�j�  j�  j  KJubK5j  )��}�(j�  K5j  ]�j�  j�  j  KJubK6j  )��}�(j�  K6j  ]�j�  j�  j  KJubK7j  )��}�(j�  K7j  ]�j�  j�  j  KJubK8j  )��}�(j�  K8j  ]�j�  j�  j  KJubK9j  )��}�(j�  K9j  ]�j�  j�  j  KJubK:j  )��}�(j�  K:j  ]�j�  j�  j  KJubK;j  )��}�(j�  K;j  ]�j�  j�  j  KJubK<j  )��}�(j�  K<j  ]�j�  j�  j  KJubK=j  )��}�(j�  K=j  ]�j�  j�  j  KJubK>j  )��}�(j�  K>j  ]�j�  j�  j  KJubK?j  )��}�(j�  K?j  ]�j�  j�  j  KJubK@j  )��}�(j�  K@j  ]�j�  j�  j  KJubKAj  )��}�(j�  KAj  ]�j�  j�  j  KJubKBj  )��}�(j�  KBj  ]�j�  j�  j  KJubKCj  )��}�(j�  KCj  ]�j�  j�  j  KJubKDj  )��}�(j�  KDj  ]�j�  j�  j  KJubKEj  )��}�(j�  KEj  ]�j�  j�  j  KJubKFj  )��}�(j�  KFj  ]�j�  j�  j  KJubKGj  )��}�(j�  KGj  ]�j�  j�  j  KJubKHj  )��}�(j�  KHj  ]�j�  j�  j  KJubKIj  )��}�(j�  KIj  ]�j�  j�  j  KJubKJj  )��}�(j�  KJj  ]�j�  j�  j  KJubKKj  )��}�(j�  KKj  ]�j�  j�  j  KJubKLj  )��}�(j�  KLj  ]�j�  j�  j  KJubKMj  )��}�(j�  KMj  ]�j�  j�  j  KJubKNj  )��}�(j�  KNj  ]�j�  j�  j  KJubKOj  )��}�(j�  KOj  ]�j�  j�  j  KJubKPj  )��}�(j�  KPj  ]�j�  j�  j  KJubKQj  )��}�(j�  KQj  ]�j�  j�  j  KJubKRj  )��}�(j�  KRj  ]�j�  j�  j  KJubKSj  )��}�(j�  KSj  ]�j�  j�  j  KJubKTj  )��}�(j�  KTj  ]�j�  j�  j  KJubKUj  )��}�(j�  KUj  ]�j�  j�  j  KJubKVj  )��}�(j�  KVj  ]�j�  j�  j  KJubKWj  )��}�(j�  KWj  ]�j�  j�  j  KJubKXj  )��}�(j�  KXj  ]�j�  j�  j  KJubKYj  )��}�(j�  KYj  ]�j�  j�  j  KJubKZj  )��}�(j�  KZj  ]�j�  j�  j  KJubK[j  )��}�(j�  K[j  ]�j�  j�  j  KJubK\j  )��}�(j�  K\j  ]�j�  j�  j  KJubK]j  )��}�(j�  K]j  ]�j�  j�  j  KJubK^j  )��}�(j�  K^j  ]�j�  j�  j  KJubK_j  )��}�(j�  K_j  ]�j�  j�  j  KJubK`j  )��}�(j�  K`j  ]�j�  j�  j  KJubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KJubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KJubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KJubuKK}�(K j  )��}�(j�  K j  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�KNaj�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�KOaj�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubK	j  )��}�(j�  K	j  ]�j�  j�  j  KKubK
j  )��}�(j�  K
j  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubKj  )��}�(j�  Kj  ]�j�  j�  j  KKubK j  )��}�(j�  K j  ]�j�  j�  j  KKubK!j  )��}�(j�  K!j  ]�j�  j�  j  KKubK"j  )��}�(j�  K"j  ]�j�  j�  j  KKubK#j  )��}�(j�  K#j  ]�j�  j�  j  KKubK$j  )��}�(j�  K$j  ]�j�  j�  j  KKubK%j  )��}�(j�  K%j  ]�j�  j�  j  KKubK&j  )��}�(j�  K&j  ]�j�  j�  j  KKubK'j  )��}�(j�  K'j  ]�j�  j�  j  KKubK(j  )��}�(j�  K(j  ]�j�  j�  j  KKubK)j  )��}�(j�  K)j  ]�j�  j�  j  KKubK*j  )��}�(j�  K*j  ]�j�  j�  j  KKubK+j  )��}�(j�  K+j  ]�j�  j�  j  KKubK,j  )��}�(j�  K,j  ]�j�  j�  j  KKubK-j  )��}�(j�  K-j  ]�j�  j�  j  KKubK.j  )��}�(j�  K.j  ]�j�  j�  j  KKubK/j  )��}�(j�  K/j  ]�j�  j�  j  KKubK0j  )��}�(j�  K0j  ]�j�  j�  j  KKubK1j  )��}�(j�  K1j  ]�j�  j�  j  KKubK2j  )��}�(j�  K2j  ]�j�  j�  j  KKubK3j  )��}�(j�  K3j  ]�j�  j�  j  KKubK4j  )��}�(j�  K4j  ]�j�  j�  j  KKubK5j  )��}�(j�  K5j  ]�j�  j�  j  KKubK6j  )��}�(j�  K6j  ]�j�  j�  j  KKubK7j  )��}�(j�  K7j  ]�j�  j�  j  KKubK8j  )��}�(j�  K8j  ]�j�  j�  j  KKubK9j  )��}�(j�  K9j  ]�j�  j�  j  KKubK:j  )��}�(j�  K:j  ]�j�  j�  j  KKubK;j  )��}�(j�  K;j  ]�j�  j�  j  KKubK<j  )��}�(j�  K<j  ]�j�  j�  j  KKubK=j  )��}�(j�  K=j  ]�j�  j�  j  KKubK>j  )��}�(j�  K>j  ]�j�  j�  j  KKubK?j  )��}�(j�  K?j  ]�j�  j�  j  KKubK@j  )��}�(j�  K@j  ]�j�  j�  j  KKubKAj  )��}�(j�  KAj  ]�j�  j�  j  KKubKBj  )��}�(j�  KBj  ]�j�  j�  j  KKubKCj  )��}�(j�  KCj  ]�j�  j�  j  KKubKDj  )��}�(j�  KDj  ]�j�  j�  j  KKubKEj  )��}�(j�  KEj  ]�j�  j�  j  KKubKFj  )��}�(j�  KFj  ]�j�  j�  j  KKubKGj  )��}�(j�  KGj  ]�j�  j�  j  KKubKHj  )��}�(j�  KHj  ]�j�  j�  j  KKubKIj  )��}�(j�  KIj  ]�j�  j�  j  KKubKJj  )��}�(j�  KJj  ]�j�  j�  j  KKubKKj  )��}�(j�  KKj  ]�j�  j�  j  KKubKLj  )��}�(j�  KLj  ]�j�  j�  j  KKubKMj  )��}�(j�  KMj  ]�j�  j�  j  KKubKNj  )��}�(j�  KNj  ]�j�  j�  j  KKubKOj  )��}�(j�  KOj  ]�j�  j�  j  KKubKPj  )��}�(j�  KPj  ]�j�  j�  j  KKubKQj  )��}�(j�  KQj  ]�j�  j�  j  KKubKRj  )��}�(j�  KRj  ]�j�  j�  j  KKubKSj  )��}�(j�  KSj  ]�j�  j�  j  KKubKTj  )��}�(j�  KTj  ]�j�  j�  j  KKubKUj  )��}�(j�  KUj  ]�j�  j�  j  KKubKVj  )��}�(j�  KVj  ]�j�  j�  j  KKubKWj  )��}�(j�  KWj  ]�j�  j�  j  KKubKXj  )��}�(j�  KXj  ]�j�  j�  j  KKubKYj  )��}�(j�  KYj  ]�j�  j�  j  KKubKZj  )��}�(j�  KZj  ]�j�  j�  j  KKubK[j  )��}�(j�  K[j  ]�j�  j�  j  KKubK\j  )��}�(j�  K\j  ]�j�  j�  j  KKubK]j  )��}�(j�  K]j  ]�j�  j�  j  KKubK^j  )��}�(j�  K^j  ]�j�  j�  j  KKubK_j  )��}�(j�  K_j  ]�j�  j�  j  KKubK`j  )��}�(j�  K`j  ]�j�  j�  j  KKubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KKubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KKubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KKubuKL}�(K j  )��}�(j�  K j  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubK	j  )��}�(j�  K	j  ]�j�  j�  j  KLubK
j  )��}�(j�  K
j  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubKj  )��}�(j�  Kj  ]�j�  j�  j  KLubK j  )��}�(j�  K j  ]�j�  j�  j  KLubK!j  )��}�(j�  K!j  ]�j�  j�  j  KLubK"j  )��}�(j�  K"j  ]�j�  j�  j  KLubK#j  )��}�(j�  K#j  ]�j�  j�  j  KLubK$j  )��}�(j�  K$j  ]�j�  j�  j  KLubK%j  )��}�(j�  K%j  ]�j�  j�  j  KLubK&j  )��}�(j�  K&j  ]�j�  j�  j  KLubK'j  )��}�(j�  K'j  ]�j�  j�  j  KLubK(j  )��}�(j�  K(j  ]�j�  j�  j  KLubK)j  )��}�(j�  K)j  ]�j�  j�  j  KLubK*j  )��}�(j�  K*j  ]�j�  j�  j  KLubK+j  )��}�(j�  K+j  ]�j�  j�  j  KLubK,j  )��}�(j�  K,j  ]�j�  j�  j  KLubK-j  )��}�(j�  K-j  ]�j�  j�  j  KLubK.j  )��}�(j�  K.j  ]�j�  j�  j  KLubK/j  )��}�(j�  K/j  ]�j�  j�  j  KLubK0j  )��}�(j�  K0j  ]�j�  j�  j  KLubK1j  )��}�(j�  K1j  ]�j�  j�  j  KLubK2j  )��}�(j�  K2j  ]�j�  j�  j  KLubK3j  )��}�(j�  K3j  ]�j�  j�  j  KLubK4j  )��}�(j�  K4j  ]�j�  j�  j  KLubK5j  )��}�(j�  K5j  ]�j�  j�  j  KLubK6j  )��}�(j�  K6j  ]�j�  j�  j  KLubK7j  )��}�(j�  K7j  ]�j�  j�  j  KLubK8j  )��}�(j�  K8j  ]�j�  j�  j  KLubK9j  )��}�(j�  K9j  ]�j�  j�  j  KLubK:j  )��}�(j�  K:j  ]�j�  j�  j  KLubK;j  )��}�(j�  K;j  ]�j�  j�  j  KLubK<j  )��}�(j�  K<j  ]�j�  j�  j  KLubK=j  )��}�(j�  K=j  ]�j�  j�  j  KLubK>j  )��}�(j�  K>j  ]�j�  j�  j  KLubK?j  )��}�(j�  K?j  ]�j�  j�  j  KLubK@j  )��}�(j�  K@j  ]�j�  j�  j  KLubKAj  )��}�(j�  KAj  ]�j�  j�  j  KLubKBj  )��}�(j�  KBj  ]�j�  j�  j  KLubKCj  )��}�(j�  KCj  ]�j�  j�  j  KLubKDj  )��}�(j�  KDj  ]�j�  j�  j  KLubKEj  )��}�(j�  KEj  ]�j�  j�  j  KLubKFj  )��}�(j�  KFj  ]�j�  j�  j  KLubKGj  )��}�(j�  KGj  ]�j�  j�  j  KLubKHj  )��}�(j�  KHj  ]�j�  j�  j  KLubKIj  )��}�(j�  KIj  ]�j�  j�  j  KLubKJj  )��}�(j�  KJj  ]�j�  j�  j  KLubKKj  )��}�(j�  KKj  ]�j�  j�  j  KLubKLj  )��}�(j�  KLj  ]�j�  j�  j  KLubKMj  )��}�(j�  KMj  ]�j�  j�  j  KLubKNj  )��}�(j�  KNj  ]�j�  j�  j  KLubKOj  )��}�(j�  KOj  ]�j�  j�  j  KLubKPj  )��}�(j�  KPj  ]�j�  j�  j  KLubKQj  )��}�(j�  KQj  ]�j�  j�  j  KLubKRj  )��}�(j�  KRj  ]�j�  j�  j  KLubKSj  )��}�(j�  KSj  ]�j�  j�  j  KLubKTj  )��}�(j�  KTj  ]�j�  j�  j  KLubKUj  )��}�(j�  KUj  ]�j�  j�  j  KLubKVj  )��}�(j�  KVj  ]�j�  j�  j  KLubKWj  )��}�(j�  KWj  ]�j�  j�  j  KLubKXj  )��}�(j�  KXj  ]�j�  j�  j  KLubKYj  )��}�(j�  KYj  ]�j�  j�  j  KLubKZj  )��}�(j�  KZj  ]�j�  j�  j  KLubK[j  )��}�(j�  K[j  ]�j�  j�  j  KLubK\j  )��}�(j�  K\j  ]�j�  j�  j  KLubK]j  )��}�(j�  K]j  ]�j�  j�  j  KLubK^j  )��}�(j�  K^j  ]�j�  j�  j  KLubK_j  )��}�(j�  K_j  ]�j�  j�  j  KLubK`j  )��}�(j�  K`j  ]�j�  j�  j  KLubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KLubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KLubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KLubuKM}�(K j  )��}�(j�  K j  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�KQaj�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubK	j  )��}�(j�  K	j  ]�j�  j�  j  KMubK
j  )��}�(j�  K
j  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubKj  )��}�(j�  Kj  ]�j�  j�  j  KMubK j  )��}�(j�  K j  ]�j�  j�  j  KMubK!j  )��}�(j�  K!j  ]�j�  j�  j  KMubK"j  )��}�(j�  K"j  ]�j�  j�  j  KMubK#j  )��}�(j�  K#j  ]�j�  j�  j  KMubK$j  )��}�(j�  K$j  ]�j�  j�  j  KMubK%j  )��}�(j�  K%j  ]�j�  j�  j  KMubK&j  )��}�(j�  K&j  ]�j�  j�  j  KMubK'j  )��}�(j�  K'j  ]�j�  j�  j  KMubK(j  )��}�(j�  K(j  ]�j�  j�  j  KMubK)j  )��}�(j�  K)j  ]�j�  j�  j  KMubK*j  )��}�(j�  K*j  ]�j�  j�  j  KMubK+j  )��}�(j�  K+j  ]�j�  j�  j  KMubK,j  )��}�(j�  K,j  ]�j�  j�  j  KMubK-j  )��}�(j�  K-j  ]�j�  j�  j  KMubK.j  )��}�(j�  K.j  ]�j�  j�  j  KMubK/j  )��}�(j�  K/j  ]�j�  j�  j  KMubK0j  )��}�(j�  K0j  ]�j�  j�  j  KMubK1j  )��}�(j�  K1j  ]�j�  j�  j  KMubK2j  )��}�(j�  K2j  ]�j�  j�  j  KMubK3j  )��}�(j�  K3j  ]�j�  j�  j  KMubK4j  )��}�(j�  K4j  ]�j�  j�  j  KMubK5j  )��}�(j�  K5j  ]�j�  j�  j  KMubK6j  )��}�(j�  K6j  ]�j�  j�  j  KMubK7j  )��}�(j�  K7j  ]�j�  j�  j  KMubK8j  )��}�(j�  K8j  ]�j�  j�  j  KMubK9j  )��}�(j�  K9j  ]�j�  j�  j  KMubK:j  )��}�(j�  K:j  ]�j�  j�  j  KMubK;j  )��}�(j�  K;j  ]�j�  j�  j  KMubK<j  )��}�(j�  K<j  ]�j�  j�  j  KMubK=j  )��}�(j�  K=j  ]�j�  j�  j  KMubK>j  )��}�(j�  K>j  ]�j�  j�  j  KMubK?j  )��}�(j�  K?j  ]�j�  j�  j  KMubK@j  )��}�(j�  K@j  ]�j�  j�  j  KMubKAj  )��}�(j�  KAj  ]�j�  j�  j  KMubKBj  )��}�(j�  KBj  ]�j�  j�  j  KMubKCj  )��}�(j�  KCj  ]�j�  j�  j  KMubKDj  )��}�(j�  KDj  ]�j�  j�  j  KMubKEj  )��}�(j�  KEj  ]�j�  j�  j  KMubKFj  )��}�(j�  KFj  ]�j�  j�  j  KMubKGj  )��}�(j�  KGj  ]�j�  j�  j  KMubKHj  )��}�(j�  KHj  ]�j�  j�  j  KMubKIj  )��}�(j�  KIj  ]�j�  j�  j  KMubKJj  )��}�(j�  KJj  ]�j�  j�  j  KMubKKj  )��}�(j�  KKj  ]�j�  j�  j  KMubKLj  )��}�(j�  KLj  ]�j�  j�  j  KMubKMj  )��}�(j�  KMj  ]�j�  j�  j  KMubKNj  )��}�(j�  KNj  ]�j�  j�  j  KMubKOj  )��}�(j�  KOj  ]�j�  j�  j  KMubKPj  )��}�(j�  KPj  ]�j�  j�  j  KMubKQj  )��}�(j�  KQj  ]�j�  j�  j  KMubKRj  )��}�(j�  KRj  ]�j�  j�  j  KMubKSj  )��}�(j�  KSj  ]�j�  j�  j  KMubKTj  )��}�(j�  KTj  ]�j�  j�  j  KMubKUj  )��}�(j�  KUj  ]�j�  j�  j  KMubKVj  )��}�(j�  KVj  ]�j�  j�  j  KMubKWj  )��}�(j�  KWj  ]�j�  j�  j  KMubKXj  )��}�(j�  KXj  ]�j�  j�  j  KMubKYj  )��}�(j�  KYj  ]�j�  j�  j  KMubKZj  )��}�(j�  KZj  ]�j�  j�  j  KMubK[j  )��}�(j�  K[j  ]�j�  j�  j  KMubK\j  )��}�(j�  K\j  ]�j�  j�  j  KMubK]j  )��}�(j�  K]j  ]�j�  j�  j  KMubK^j  )��}�(j�  K^j  ]�j�  j�  j  KMubK_j  )��}�(j�  K_j  ]�j�  j�  j  KMubK`j  )��}�(j�  K`j  ]�j�  j�  j  KMubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KMubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KMubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KMubuKN}�(K j  )��}�(j�  K j  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�KRaj�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�KSaj�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubK	j  )��}�(j�  K	j  ]�j�  j�  j  KNubK
j  )��}�(j�  K
j  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubKj  )��}�(j�  Kj  ]�j�  j�  j  KNubK j  )��}�(j�  K j  ]�j�  j�  j  KNubK!j  )��}�(j�  K!j  ]�j�  j�  j  KNubK"j  )��}�(j�  K"j  ]�j�  j�  j  KNubK#j  )��}�(j�  K#j  ]�j�  j�  j  KNubK$j  )��}�(j�  K$j  ]�j�  j�  j  KNubK%j  )��}�(j�  K%j  ]�j�  j�  j  KNubK&j  )��}�(j�  K&j  ]�j�  j�  j  KNubK'j  )��}�(j�  K'j  ]�j�  j�  j  KNubK(j  )��}�(j�  K(j  ]�j�  j�  j  KNubK)j  )��}�(j�  K)j  ]�j�  j�  j  KNubK*j  )��}�(j�  K*j  ]�j�  j�  j  KNubK+j  )��}�(j�  K+j  ]�j�  j�  j  KNubK,j  )��}�(j�  K,j  ]�j�  j�  j  KNubK-j  )��}�(j�  K-j  ]�j�  j�  j  KNubK.j  )��}�(j�  K.j  ]�j�  j�  j  KNubK/j  )��}�(j�  K/j  ]�j�  j�  j  KNubK0j  )��}�(j�  K0j  ]�j�  j�  j  KNubK1j  )��}�(j�  K1j  ]�j�  j�  j  KNubK2j  )��}�(j�  K2j  ]�j�  j�  j  KNubK3j  )��}�(j�  K3j  ]�j�  j�  j  KNubK4j  )��}�(j�  K4j  ]�j�  j�  j  KNubK5j  )��}�(j�  K5j  ]�j�  j�  j  KNubK6j  )��}�(j�  K6j  ]�j�  j�  j  KNubK7j  )��}�(j�  K7j  ]�j�  j�  j  KNubK8j  )��}�(j�  K8j  ]�j�  j�  j  KNubK9j  )��}�(j�  K9j  ]�j�  j�  j  KNubK:j  )��}�(j�  K:j  ]�j�  j�  j  KNubK;j  )��}�(j�  K;j  ]�j�  j�  j  KNubK<j  )��}�(j�  K<j  ]�j�  j�  j  KNubK=j  )��}�(j�  K=j  ]�j�  j�  j  KNubK>j  )��}�(j�  K>j  ]�j�  j�  j  KNubK?j  )��}�(j�  K?j  ]�j�  j�  j  KNubK@j  )��}�(j�  K@j  ]�j�  j�  j  KNubKAj  )��}�(j�  KAj  ]�j�  j�  j  KNubKBj  )��}�(j�  KBj  ]�j�  j�  j  KNubKCj  )��}�(j�  KCj  ]�j�  j�  j  KNubKDj  )��}�(j�  KDj  ]�j�  j�  j  KNubKEj  )��}�(j�  KEj  ]�j�  j�  j  KNubKFj  )��}�(j�  KFj  ]�j�  j�  j  KNubKGj  )��}�(j�  KGj  ]�j�  j�  j  KNubKHj  )��}�(j�  KHj  ]�j�  j�  j  KNubKIj  )��}�(j�  KIj  ]�j�  j�  j  KNubKJj  )��}�(j�  KJj  ]�j�  j�  j  KNubKKj  )��}�(j�  KKj  ]�j�  j�  j  KNubKLj  )��}�(j�  KLj  ]�j�  j�  j  KNubKMj  )��}�(j�  KMj  ]�j�  j�  j  KNubKNj  )��}�(j�  KNj  ]�j�  j�  j  KNubKOj  )��}�(j�  KOj  ]�j�  j�  j  KNubKPj  )��}�(j�  KPj  ]�j�  j�  j  KNubKQj  )��}�(j�  KQj  ]�j�  j�  j  KNubKRj  )��}�(j�  KRj  ]�j�  j�  j  KNubKSj  )��}�(j�  KSj  ]�j�  j�  j  KNubKTj  )��}�(j�  KTj  ]�j�  j�  j  KNubKUj  )��}�(j�  KUj  ]�j�  j�  j  KNubKVj  )��}�(j�  KVj  ]�j�  j�  j  KNubKWj  )��}�(j�  KWj  ]�j�  j�  j  KNubKXj  )��}�(j�  KXj  ]�j�  j�  j  KNubKYj  )��}�(j�  KYj  ]�j�  j�  j  KNubKZj  )��}�(j�  KZj  ]�j�  j�  j  KNubK[j  )��}�(j�  K[j  ]�j�  j�  j  KNubK\j  )��}�(j�  K\j  ]�j�  j�  j  KNubK]j  )��}�(j�  K]j  ]�j�  j�  j  KNubK^j  )��}�(j�  K^j  ]�j�  j�  j  KNubK_j  )��}�(j�  K_j  ]�j�  j�  j  KNubK`j  )��}�(j�  K`j  ]�j�  j�  j  KNubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KNubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KNubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KNubuKO}�(K j  )��}�(j�  K j  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubK	j  )��}�(j�  K	j  ]�j�  j�  j  KOubK
j  )��}�(j�  K
j  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�KTaj�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubKj  )��}�(j�  Kj  ]�j�  j�  j  KOubK j  )��}�(j�  K j  ]�j�  j�  j  KOubK!j  )��}�(j�  K!j  ]�j�  j�  j  KOubK"j  )��}�(j�  K"j  ]�j�  j�  j  KOubK#j  )��}�(j�  K#j  ]�j�  j�  j  KOubK$j  )��}�(j�  K$j  ]�j�  j�  j  KOubK%j  )��}�(j�  K%j  ]�j�  j�  j  KOubK&j  )��}�(j�  K&j  ]�j�  j�  j  KOubK'j  )��}�(j�  K'j  ]�j�  j�  j  KOubK(j  )��}�(j�  K(j  ]�j�  j�  j  KOubK)j  )��}�(j�  K)j  ]�j�  j�  j  KOubK*j  )��}�(j�  K*j  ]�j�  j�  j  KOubK+j  )��}�(j�  K+j  ]�j�  j�  j  KOubK,j  )��}�(j�  K,j  ]�j�  j�  j  KOubK-j  )��}�(j�  K-j  ]�j�  j�  j  KOubK.j  )��}�(j�  K.j  ]�j�  j�  j  KOubK/j  )��}�(j�  K/j  ]�j�  j�  j  KOubK0j  )��}�(j�  K0j  ]�j�  j�  j  KOubK1j  )��}�(j�  K1j  ]�j�  j�  j  KOubK2j  )��}�(j�  K2j  ]�j�  j�  j  KOubK3j  )��}�(j�  K3j  ]�j�  j�  j  KOubK4j  )��}�(j�  K4j  ]�j�  j�  j  KOubK5j  )��}�(j�  K5j  ]�j�  j�  j  KOubK6j  )��}�(j�  K6j  ]�j�  j�  j  KOubK7j  )��}�(j�  K7j  ]�j�  j�  j  KOubK8j  )��}�(j�  K8j  ]�j�  j�  j  KOubK9j  )��}�(j�  K9j  ]�j�  j�  j  KOubK:j  )��}�(j�  K:j  ]�j�  j�  j  KOubK;j  )��}�(j�  K;j  ]�j�  j�  j  KOubK<j  )��}�(j�  K<j  ]�j�  j�  j  KOubK=j  )��}�(j�  K=j  ]�j�  j�  j  KOubK>j  )��}�(j�  K>j  ]�j�  j�  j  KOubK?j  )��}�(j�  K?j  ]�j�  j�  j  KOubK@j  )��}�(j�  K@j  ]�j�  j�  j  KOubKAj  )��}�(j�  KAj  ]�j�  j�  j  KOubKBj  )��}�(j�  KBj  ]�j�  j�  j  KOubKCj  )��}�(j�  KCj  ]�j�  j�  j  KOubKDj  )��}�(j�  KDj  ]�j�  j�  j  KOubKEj  )��}�(j�  KEj  ]�j�  j�  j  KOubKFj  )��}�(j�  KFj  ]�j�  j�  j  KOubKGj  )��}�(j�  KGj  ]�j�  j�  j  KOubKHj  )��}�(j�  KHj  ]�j�  j�  j  KOubKIj  )��}�(j�  KIj  ]�j�  j�  j  KOubKJj  )��}�(j�  KJj  ]�j�  j�  j  KOubKKj  )��}�(j�  KKj  ]�j�  j�  j  KOubKLj  )��}�(j�  KLj  ]�KVaj�  j�  j  KOubKMj  )��}�(j�  KMj  ]�j�  j�  j  KOubKNj  )��}�(j�  KNj  ]�j�  j�  j  KOubKOj  )��}�(j�  KOj  ]�j�  j�  j  KOubKPj  )��}�(j�  KPj  ]�j�  j�  j  KOubKQj  )��}�(j�  KQj  ]�j�  j�  j  KOubKRj  )��}�(j�  KRj  ]�j�  j�  j  KOubKSj  )��}�(j�  KSj  ]�j�  j�  j  KOubKTj  )��}�(j�  KTj  ]�j�  j�  j  KOubKUj  )��}�(j�  KUj  ]�j�  j�  j  KOubKVj  )��}�(j�  KVj  ]�j�  j�  j  KOubKWj  )��}�(j�  KWj  ]�j�  j�  j  KOubKXj  )��}�(j�  KXj  ]�j�  j�  j  KOubKYj  )��}�(j�  KYj  ]�j�  j�  j  KOubKZj  )��}�(j�  KZj  ]�j�  j�  j  KOubK[j  )��}�(j�  K[j  ]�j�  j�  j  KOubK\j  )��}�(j�  K\j  ]�j�  j�  j  KOubK]j  )��}�(j�  K]j  ]�j�  j�  j  KOubK^j  )��}�(j�  K^j  ]�j�  j�  j  KOubK_j  )��}�(j�  K_j  ]�j�  j�  j  KOubK`j  )��}�(j�  K`j  ]�j�  j�  j  KOubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KOubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KOubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KOubuKP}�(K j  )��}�(j�  K j  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubK	j  )��}�(j�  K	j  ]�j�  j�  j  KPubK
j  )��}�(j�  K
j  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�KXaj�  j�  j  KPubKj  )��}�(j�  Kj  ]�KYaj�  j�  j  KPubKj  )��}�(j�  Kj  ]�KZaj�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubKj  )��}�(j�  Kj  ]�j�  j�  j  KPubK j  )��}�(j�  K j  ]�j�  j�  j  KPubK!j  )��}�(j�  K!j  ]�j�  j�  j  KPubK"j  )��}�(j�  K"j  ]�j�  j�  j  KPubK#j  )��}�(j�  K#j  ]�j�  j�  j  KPubK$j  )��}�(j�  K$j  ]�j�  j�  j  KPubK%j  )��}�(j�  K%j  ]�j�  j�  j  KPubK&j  )��}�(j�  K&j  ]�j�  j�  j  KPubK'j  )��}�(j�  K'j  ]�j�  j�  j  KPubK(j  )��}�(j�  K(j  ]�j�  j�  j  KPubK)j  )��}�(j�  K)j  ]�j�  j�  j  KPubK*j  )��}�(j�  K*j  ]�j�  j�  j  KPubK+j  )��}�(j�  K+j  ]�j�  j�  j  KPubK,j  )��}�(j�  K,j  ]�j�  j�  j  KPubK-j  )��}�(j�  K-j  ]�j�  j�  j  KPubK.j  )��}�(j�  K.j  ]�j�  j�  j  KPubK/j  )��}�(j�  K/j  ]�j�  j�  j  KPubK0j  )��}�(j�  K0j  ]�j�  j�  j  KPubK1j  )��}�(j�  K1j  ]�j�  j�  j  KPubK2j  )��}�(j�  K2j  ]�j�  j�  j  KPubK3j  )��}�(j�  K3j  ]�j�  j�  j  KPubK4j  )��}�(j�  K4j  ]�j�  j�  j  KPubK5j  )��}�(j�  K5j  ]�j�  j�  j  KPubK6j  )��}�(j�  K6j  ]�j�  j�  j  KPubK7j  )��}�(j�  K7j  ]�j�  j�  j  KPubK8j  )��}�(j�  K8j  ]�j�  j�  j  KPubK9j  )��}�(j�  K9j  ]�j�  j�  j  KPubK:j  )��}�(j�  K:j  ]�j�  j�  j  KPubK;j  )��}�(j�  K;j  ]�j�  j�  j  KPubK<j  )��}�(j�  K<j  ]�j�  j�  j  KPubK=j  )��}�(j�  K=j  ]�j�  j�  j  KPubK>j  )��}�(j�  K>j  ]�j�  j�  j  KPubK?j  )��}�(j�  K?j  ]�j�  j�  j  KPubK@j  )��}�(j�  K@j  ]�j�  j�  j  KPubKAj  )��}�(j�  KAj  ]�j�  j�  j  KPubKBj  )��}�(j�  KBj  ]�j�  j�  j  KPubKCj  )��}�(j�  KCj  ]�j�  j�  j  KPubKDj  )��}�(j�  KDj  ]�j�  j�  j  KPubKEj  )��}�(j�  KEj  ]�j�  j�  j  KPubKFj  )��}�(j�  KFj  ]�j�  j�  j  KPubKGj  )��}�(j�  KGj  ]�j�  j�  j  KPubKHj  )��}�(j�  KHj  ]�j�  j�  j  KPubKIj  )��}�(j�  KIj  ]�j�  j�  j  KPubKJj  )��}�(j�  KJj  ]�j�  j�  j  KPubKKj  )��}�(j�  KKj  ]�j�  j�  j  KPubKLj  )��}�(j�  KLj  ]�j�  j�  j  KPubKMj  )��}�(j�  KMj  ]�j�  j�  j  KPubKNj  )��}�(j�  KNj  ]�j�  j�  j  KPubKOj  )��}�(j�  KOj  ]�j�  j�  j  KPubKPj  )��}�(j�  KPj  ]�j�  j�  j  KPubKQj  )��}�(j�  KQj  ]�j�  j�  j  KPubKRj  )��}�(j�  KRj  ]�j�  j�  j  KPubKSj  )��}�(j�  KSj  ]�j�  j�  j  KPubKTj  )��}�(j�  KTj  ]�j�  j�  j  KPubKUj  )��}�(j�  KUj  ]�j�  j�  j  KPubKVj  )��}�(j�  KVj  ]�j�  j�  j  KPubKWj  )��}�(j�  KWj  ]�j�  j�  j  KPubKXj  )��}�(j�  KXj  ]�j�  j�  j  KPubKYj  )��}�(j�  KYj  ]�j�  j�  j  KPubKZj  )��}�(j�  KZj  ]�j�  j�  j  KPubK[j  )��}�(j�  K[j  ]�j�  j�  j  KPubK\j  )��}�(j�  K\j  ]�j�  j�  j  KPubK]j  )��}�(j�  K]j  ]�j�  j�  j  KPubK^j  )��}�(j�  K^j  ]�j�  j�  j  KPubK_j  )��}�(j�  K_j  ]�j�  j�  j  KPubK`j  )��}�(j�  K`j  ]�j�  j�  j  KPubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KPubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KPubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KPubuKQ}�(K j  )��}�(j�  K j  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubK	j  )��}�(j�  K	j  ]�j�  j�  j  KQubK
j  )��}�(j�  K
j  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�K]aj�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubKj  )��}�(j�  Kj  ]�j�  j�  j  KQubK j  )��}�(j�  K j  ]�j�  j�  j  KQubK!j  )��}�(j�  K!j  ]�j�  j�  j  KQubK"j  )��}�(j�  K"j  ]�j�  j�  j  KQubK#j  )��}�(j�  K#j  ]�j�  j�  j  KQubK$j  )��}�(j�  K$j  ]�j�  j�  j  KQubK%j  )��}�(j�  K%j  ]�j�  j�  j  KQubK&j  )��}�(j�  K&j  ]�j�  j�  j  KQubK'j  )��}�(j�  K'j  ]�j�  j�  j  KQubK(j  )��}�(j�  K(j  ]�j�  j�  j  KQubK)j  )��}�(j�  K)j  ]�j�  j�  j  KQubK*j  )��}�(j�  K*j  ]�j�  j�  j  KQubK+j  )��}�(j�  K+j  ]�j�  j�  j  KQubK,j  )��}�(j�  K,j  ]�j�  j�  j  KQubK-j  )��}�(j�  K-j  ]�j�  j�  j  KQubK.j  )��}�(j�  K.j  ]�j�  j�  j  KQubK/j  )��}�(j�  K/j  ]�j�  j�  j  KQubK0j  )��}�(j�  K0j  ]�j�  j�  j  KQubK1j  )��}�(j�  K1j  ]�j�  j�  j  KQubK2j  )��}�(j�  K2j  ]�j�  j�  j  KQubK3j  )��}�(j�  K3j  ]�j�  j�  j  KQubK4j  )��}�(j�  K4j  ]�j�  j�  j  KQubK5j  )��}�(j�  K5j  ]�j�  j�  j  KQubK6j  )��}�(j�  K6j  ]�j�  j�  j  KQubK7j  )��}�(j�  K7j  ]�j�  j�  j  KQubK8j  )��}�(j�  K8j  ]�j�  j�  j  KQubK9j  )��}�(j�  K9j  ]�j�  j�  j  KQubK:j  )��}�(j�  K:j  ]�j�  j�  j  KQubK;j  )��}�(j�  K;j  ]�j�  j�  j  KQubK<j  )��}�(j�  K<j  ]�j�  j�  j  KQubK=j  )��}�(j�  K=j  ]�j�  j�  j  KQubK>j  )��}�(j�  K>j  ]�j�  j�  j  KQubK?j  )��}�(j�  K?j  ]�j�  j�  j  KQubK@j  )��}�(j�  K@j  ]�j�  j�  j  KQubKAj  )��}�(j�  KAj  ]�j�  j�  j  KQubKBj  )��}�(j�  KBj  ]�j�  j�  j  KQubKCj  )��}�(j�  KCj  ]�j�  j�  j  KQubKDj  )��}�(j�  KDj  ]�j�  j�  j  KQubKEj  )��}�(j�  KEj  ]�j�  j�  j  KQubKFj  )��}�(j�  KFj  ]�j�  j�  j  KQubKGj  )��}�(j�  KGj  ]�j�  j�  j  KQubKHj  )��}�(j�  KHj  ]�j�  j�  j  KQubKIj  )��}�(j�  KIj  ]�j�  j�  j  KQubKJj  )��}�(j�  KJj  ]�j�  j�  j  KQubKKj  )��}�(j�  KKj  ]�j�  j�  j  KQubKLj  )��}�(j�  KLj  ]�j�  j�  j  KQubKMj  )��}�(j�  KMj  ]�j�  j�  j  KQubKNj  )��}�(j�  KNj  ]�j�  j�  j  KQubKOj  )��}�(j�  KOj  ]�j�  j�  j  KQubKPj  )��}�(j�  KPj  ]�j�  j�  j  KQubKQj  )��}�(j�  KQj  ]�j�  j�  j  KQubKRj  )��}�(j�  KRj  ]�j�  j�  j  KQubKSj  )��}�(j�  KSj  ]�j�  j�  j  KQubKTj  )��}�(j�  KTj  ]�j�  j�  j  KQubKUj  )��}�(j�  KUj  ]�j�  j�  j  KQubKVj  )��}�(j�  KVj  ]�j�  j�  j  KQubKWj  )��}�(j�  KWj  ]�j�  j�  j  KQubKXj  )��}�(j�  KXj  ]�j�  j�  j  KQubKYj  )��}�(j�  KYj  ]�j�  j�  j  KQubKZj  )��}�(j�  KZj  ]�j�  j�  j  KQubK[j  )��}�(j�  K[j  ]�j�  j�  j  KQubK\j  )��}�(j�  K\j  ]�j�  j�  j  KQubK]j  )��}�(j�  K]j  ]�j�  j�  j  KQubK^j  )��}�(j�  K^j  ]�j�  j�  j  KQubK_j  )��}�(j�  K_j  ]�j�  j�  j  KQubK`j  )��}�(j�  K`j  ]�j�  j�  j  KQubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KQubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KQubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KQubuKR}�(K j  )��}�(j�  K j  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubK	j  )��}�(j�  K	j  ]�j�  j�  j  KRubK
j  )��}�(j�  K
j  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�Kbaj�  j�  j  KRubKj  )��}�(j�  Kj  ]�Kcaj�  j�  j  KRubKj  )��}�(j�  Kj  ]�Kdaj�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubKj  )��}�(j�  Kj  ]�j�  j�  j  KRubK j  )��}�(j�  K j  ]�j�  j�  j  KRubK!j  )��}�(j�  K!j  ]�j�  j�  j  KRubK"j  )��}�(j�  K"j  ]�j�  j�  j  KRubK#j  )��}�(j�  K#j  ]�j�  j�  j  KRubK$j  )��}�(j�  K$j  ]�j�  j�  j  KRubK%j  )��}�(j�  K%j  ]�j�  j�  j  KRubK&j  )��}�(j�  K&j  ]�j�  j�  j  KRubK'j  )��}�(j�  K'j  ]�j�  j�  j  KRubK(j  )��}�(j�  K(j  ]�j�  j�  j  KRubK)j  )��}�(j�  K)j  ]�j�  j�  j  KRubK*j  )��}�(j�  K*j  ]�j�  j�  j  KRubK+j  )��}�(j�  K+j  ]�j�  j�  j  KRubK,j  )��}�(j�  K,j  ]�j�  j�  j  KRubK-j  )��}�(j�  K-j  ]�j�  j�  j  KRubK.j  )��}�(j�  K.j  ]�j�  j�  j  KRubK/j  )��}�(j�  K/j  ]�j�  j�  j  KRubK0j  )��}�(j�  K0j  ]�j�  j�  j  KRubK1j  )��}�(j�  K1j  ]�j�  j�  j  KRubK2j  )��}�(j�  K2j  ]�j�  j�  j  KRubK3j  )��}�(j�  K3j  ]�j�  j�  j  KRubK4j  )��}�(j�  K4j  ]�j�  j�  j  KRubK5j  )��}�(j�  K5j  ]�j�  j�  j  KRubK6j  )��}�(j�  K6j  ]�j�  j�  j  KRubK7j  )��}�(j�  K7j  ]�j�  j�  j  KRubK8j  )��}�(j�  K8j  ]�j�  j�  j  KRubK9j  )��}�(j�  K9j  ]�j�  j�  j  KRubK:j  )��}�(j�  K:j  ]�j�  j�  j  KRubK;j  )��}�(j�  K;j  ]�j�  j�  j  KRubK<j  )��}�(j�  K<j  ]�j�  j�  j  KRubK=j  )��}�(j�  K=j  ]�j�  j�  j  KRubK>j  )��}�(j�  K>j  ]�j�  j�  j  KRubK?j  )��}�(j�  K?j  ]�j�  j�  j  KRubK@j  )��}�(j�  K@j  ]�j�  j�  j  KRubKAj  )��}�(j�  KAj  ]�j�  j�  j  KRubKBj  )��}�(j�  KBj  ]�j�  j�  j  KRubKCj  )��}�(j�  KCj  ]�(K�K�ej�  j�  j  KRubKDj  )��}�(j�  KDj  ]�j�  j�  j  KRubKEj  )��}�(j�  KEj  ]�KFaj�  j�  j  KRubKFj  )��}�(j�  KFj  ]�(K�K�K�ej�  j�  j  KRubKGj  )��}�(j�  KGj  ]�j�  j�  j  KRubKHj  )��}�(j�  KHj  ]�j�  j�  j  KRubKIj  )��}�(j�  KIj  ]�j�  j�  j  KRubKJj  )��}�(j�  KJj  ]�j�  j�  j  KRubKKj  )��}�(j�  KKj  ]�j�  j�  j  KRubKLj  )��}�(j�  KLj  ]�j�  j�  j  KRubKMj  )��}�(j�  KMj  ]�j�  j�  j  KRubKNj  )��}�(j�  KNj  ]�j�  j�  j  KRubKOj  )��}�(j�  KOj  ]�j�  j�  j  KRubKPj  )��}�(j�  KPj  ]�j�  j�  j  KRubKQj  )��}�(j�  KQj  ]�j�  j�  j  KRubKRj  )��}�(j�  KRj  ]�j�  j�  j  KRubKSj  )��}�(j�  KSj  ]�j�  j�  j  KRubKTj  )��}�(j�  KTj  ]�j�  j�  j  KRubKUj  )��}�(j�  KUj  ]�j�  j�  j  KRubKVj  )��}�(j�  KVj  ]�j�  j�  j  KRubKWj  )��}�(j�  KWj  ]�j�  j�  j  KRubKXj  )��}�(j�  KXj  ]�j�  j�  j  KRubKYj  )��}�(j�  KYj  ]�j�  j�  j  KRubKZj  )��}�(j�  KZj  ]�j�  j�  j  KRubK[j  )��}�(j�  K[j  ]�j�  j�  j  KRubK\j  )��}�(j�  K\j  ]�j�  j�  j  KRubK]j  )��}�(j�  K]j  ]�j�  j�  j  KRubK^j  )��}�(j�  K^j  ]�j�  j�  j  KRubK_j  )��}�(j�  K_j  ]�j�  j�  j  KRubK`j  )��}�(j�  K`j  ]�j�  j�  j  KRubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KRubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KRubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KRubuKS}�(K j  )��}�(j�  K j  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubK	j  )��}�(j�  K	j  ]�j�  j�  j  KSubK
j  )��}�(j�  K
j  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubKj  )��}�(j�  Kj  ]�j�  j�  j  KSubK j  )��}�(j�  K j  ]�j�  j�  j  KSubK!j  )��}�(j�  K!j  ]�j�  j�  j  KSubK"j  )��}�(j�  K"j  ]�j�  j�  j  KSubK#j  )��}�(j�  K#j  ]�j�  j�  j  KSubK$j  )��}�(j�  K$j  ]�j�  j�  j  KSubK%j  )��}�(j�  K%j  ]�j�  j�  j  KSubK&j  )��}�(j�  K&j  ]�j�  j�  j  KSubK'j  )��}�(j�  K'j  ]�j�  j�  j  KSubK(j  )��}�(j�  K(j  ]�j�  j�  j  KSubK)j  )��}�(j�  K)j  ]�j�  j�  j  KSubK*j  )��}�(j�  K*j  ]�j�  j�  j  KSubK+j  )��}�(j�  K+j  ]�j�  j�  j  KSubK,j  )��}�(j�  K,j  ]�j�  j�  j  KSubK-j  )��}�(j�  K-j  ]�j�  j�  j  KSubK.j  )��}�(j�  K.j  ]�j�  j�  j  KSubK/j  )��}�(j�  K/j  ]�j�  j�  j  KSubK0j  )��}�(j�  K0j  ]�j�  j�  j  KSubK1j  )��}�(j�  K1j  ]�j�  j�  j  KSubK2j  )��}�(j�  K2j  ]�j�  j�  j  KSubK3j  )��}�(j�  K3j  ]�j�  j�  j  KSubK4j  )��}�(j�  K4j  ]�j�  j�  j  KSubK5j  )��}�(j�  K5j  ]�j�  j�  j  KSubK6j  )��}�(j�  K6j  ]�j�  j�  j  KSubK7j  )��}�(j�  K7j  ]�j�  j�  j  KSubK8j  )��}�(j�  K8j  ]�j�  j�  j  KSubK9j  )��}�(j�  K9j  ]�j�  j�  j  KSubK:j  )��}�(j�  K:j  ]�j�  j�  j  KSubK;j  )��}�(j�  K;j  ]�j�  j�  j  KSubK<j  )��}�(j�  K<j  ]�j�  j�  j  KSubK=j  )��}�(j�  K=j  ]�j�  j�  j  KSubK>j  )��}�(j�  K>j  ]�j�  j�  j  KSubK?j  )��}�(j�  K?j  ]�j�  j�  j  KSubK@j  )��}�(j�  K@j  ]�j�  j�  j  KSubKAj  )��}�(j�  KAj  ]�j�  j�  j  KSubKBj  )��}�(j�  KBj  ]�j�  j�  j  KSubKCj  )��}�(j�  KCj  ]�j�  j�  j  KSubKDj  )��}�(j�  KDj  ]�j�  j�  j  KSubKEj  )��}�(j�  KEj  ]�j�  j�  j  KSubKFj  )��}�(j�  KFj  ]�j�  j�  j  KSubKGj  )��}�(j�  KGj  ]�j�  j�  j  KSubKHj  )��}�(j�  KHj  ]�j�  j�  j  KSubKIj  )��}�(j�  KIj  ]�j�  j�  j  KSubKJj  )��}�(j�  KJj  ]�j�  j�  j  KSubKKj  )��}�(j�  KKj  ]�j�  j�  j  KSubKLj  )��}�(j�  KLj  ]�j�  j�  j  KSubKMj  )��}�(j�  KMj  ]�j�  j�  j  KSubKNj  )��}�(j�  KNj  ]�j�  j�  j  KSubKOj  )��}�(j�  KOj  ]�Khaj�  j�  j  KSubKPj  )��}�(j�  KPj  ]�j�  j�  j  KSubKQj  )��}�(j�  KQj  ]�j�  j�  j  KSubKRj  )��}�(j�  KRj  ]�j�  j�  j  KSubKSj  )��}�(j�  KSj  ]�j�  j�  j  KSubKTj  )��}�(j�  KTj  ]�j�  j�  j  KSubKUj  )��}�(j�  KUj  ]�j�  j�  j  KSubKVj  )��}�(j�  KVj  ]�j�  j�  j  KSubKWj  )��}�(j�  KWj  ]�j�  j�  j  KSubKXj  )��}�(j�  KXj  ]�j�  j�  j  KSubKYj  )��}�(j�  KYj  ]�j�  j�  j  KSubKZj  )��}�(j�  KZj  ]�j�  j�  j  KSubK[j  )��}�(j�  K[j  ]�j�  j�  j  KSubK\j  )��}�(j�  K\j  ]�j�  j�  j  KSubK]j  )��}�(j�  K]j  ]�j�  j�  j  KSubK^j  )��}�(j�  K^j  ]�j�  j�  j  KSubK_j  )��}�(j�  K_j  ]�j�  j�  j  KSubK`j  )��}�(j�  K`j  ]�j�  j�  j  KSubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KSubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KSubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KSubuKT}�(K j  )��}�(j�  K j  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubK	j  )��}�(j�  K	j  ]�j�  j�  j  KTubK
j  )��}�(j�  K
j  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubKj  )��}�(j�  Kj  ]�j�  j�  j  KTubK j  )��}�(j�  K j  ]�j�  j�  j  KTubK!j  )��}�(j�  K!j  ]�j�  j�  j  KTubK"j  )��}�(j�  K"j  ]�j�  j�  j  KTubK#j  )��}�(j�  K#j  ]�j�  j�  j  KTubK$j  )��}�(j�  K$j  ]�j�  j�  j  KTubK%j  )��}�(j�  K%j  ]�j�  j�  j  KTubK&j  )��}�(j�  K&j  ]�j�  j�  j  KTubK'j  )��}�(j�  K'j  ]�j�  j�  j  KTubK(j  )��}�(j�  K(j  ]�j�  j�  j  KTubK)j  )��}�(j�  K)j  ]�j�  j�  j  KTubK*j  )��}�(j�  K*j  ]�j�  j�  j  KTubK+j  )��}�(j�  K+j  ]�j�  j�  j  KTubK,j  )��}�(j�  K,j  ]�j�  j�  j  KTubK-j  )��}�(j�  K-j  ]�j�  j�  j  KTubK.j  )��}�(j�  K.j  ]�j�  j�  j  KTubK/j  )��}�(j�  K/j  ]�j�  j�  j  KTubK0j  )��}�(j�  K0j  ]�j�  j�  j  KTubK1j  )��}�(j�  K1j  ]�j�  j�  j  KTubK2j  )��}�(j�  K2j  ]�j�  j�  j  KTubK3j  )��}�(j�  K3j  ]�j�  j�  j  KTubK4j  )��}�(j�  K4j  ]�j�  j�  j  KTubK5j  )��}�(j�  K5j  ]�j�  j�  j  KTubK6j  )��}�(j�  K6j  ]�j�  j�  j  KTubK7j  )��}�(j�  K7j  ]�j�  j�  j  KTubK8j  )��}�(j�  K8j  ]�j�  j�  j  KTubK9j  )��}�(j�  K9j  ]�j�  j�  j  KTubK:j  )��}�(j�  K:j  ]�j�  j�  j  KTubK;j  )��}�(j�  K;j  ]�j�  j�  j  KTubK<j  )��}�(j�  K<j  ]�j�  j�  j  KTubK=j  )��}�(j�  K=j  ]�j�  j�  j  KTubK>j  )��}�(j�  K>j  ]�j�  j�  j  KTubK?j  )��}�(j�  K?j  ]�j�  j�  j  KTubK@j  )��}�(j�  K@j  ]�j�  j�  j  KTubKAj  )��}�(j�  KAj  ]�j�  j�  j  KTubKBj  )��}�(j�  KBj  ]�j�  j�  j  KTubKCj  )��}�(j�  KCj  ]�j�  j�  j  KTubKDj  )��}�(j�  KDj  ]�j�  j�  j  KTubKEj  )��}�(j�  KEj  ]�j�  j�  j  KTubKFj  )��}�(j�  KFj  ]�j�  j�  j  KTubKGj  )��}�(j�  KGj  ]�j�  j�  j  KTubKHj  )��}�(j�  KHj  ]�j�  j�  j  KTubKIj  )��}�(j�  KIj  ]�j�  j�  j  KTubKJj  )��}�(j�  KJj  ]�j�  j�  j  KTubKKj  )��}�(j�  KKj  ]�j�  j�  j  KTubKLj  )��}�(j�  KLj  ]�j�  j�  j  KTubKMj  )��}�(j�  KMj  ]�j�  j�  j  KTubKNj  )��}�(j�  KNj  ]�j�  j�  j  KTubKOj  )��}�(j�  KOj  ]�j�  j�  j  KTubKPj  )��}�(j�  KPj  ]�j�  j�  j  KTubKQj  )��}�(j�  KQj  ]�j�  j�  j  KTubKRj  )��}�(j�  KRj  ]�j�  j�  j  KTubKSj  )��}�(j�  KSj  ]�j�  j�  j  KTubKTj  )��}�(j�  KTj  ]�j�  j�  j  KTubKUj  )��}�(j�  KUj  ]�j�  j�  j  KTubKVj  )��}�(j�  KVj  ]�j�  j�  j  KTubKWj  )��}�(j�  KWj  ]�j�  j�  j  KTubKXj  )��}�(j�  KXj  ]�j�  j�  j  KTubKYj  )��}�(j�  KYj  ]�j�  j�  j  KTubKZj  )��}�(j�  KZj  ]�j�  j�  j  KTubK[j  )��}�(j�  K[j  ]�j�  j�  j  KTubK\j  )��}�(j�  K\j  ]�j�  j�  j  KTubK]j  )��}�(j�  K]j  ]�j�  j�  j  KTubK^j  )��}�(j�  K^j  ]�j�  j�  j  KTubK_j  )��}�(j�  K_j  ]�j�  j�  j  KTubK`j  )��}�(j�  K`j  ]�j�  j�  j  KTubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KTubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KTubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KTubuKU}�(K j  )��}�(j�  K j  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubK	j  )��}�(j�  K	j  ]�j�  j�  j  KUubK
j  )��}�(j�  K
j  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubKj  )��}�(j�  Kj  ]�j�  j�  j  KUubK j  )��}�(j�  K j  ]�j�  j�  j  KUubK!j  )��}�(j�  K!j  ]�j�  j�  j  KUubK"j  )��}�(j�  K"j  ]�j�  j�  j  KUubK#j  )��}�(j�  K#j  ]�j�  j�  j  KUubK$j  )��}�(j�  K$j  ]�j�  j�  j  KUubK%j  )��}�(j�  K%j  ]�j�  j�  j  KUubK&j  )��}�(j�  K&j  ]�j�  j�  j  KUubK'j  )��}�(j�  K'j  ]�j�  j�  j  KUubK(j  )��}�(j�  K(j  ]�j�  j�  j  KUubK)j  )��}�(j�  K)j  ]�j�  j�  j  KUubK*j  )��}�(j�  K*j  ]�j�  j�  j  KUubK+j  )��}�(j�  K+j  ]�j�  j�  j  KUubK,j  )��}�(j�  K,j  ]�j�  j�  j  KUubK-j  )��}�(j�  K-j  ]�j�  j�  j  KUubK.j  )��}�(j�  K.j  ]�j�  j�  j  KUubK/j  )��}�(j�  K/j  ]�j�  j�  j  KUubK0j  )��}�(j�  K0j  ]�j�  j�  j  KUubK1j  )��}�(j�  K1j  ]�j�  j�  j  KUubK2j  )��}�(j�  K2j  ]�j�  j�  j  KUubK3j  )��}�(j�  K3j  ]�j�  j�  j  KUubK4j  )��}�(j�  K4j  ]�j�  j�  j  KUubK5j  )��}�(j�  K5j  ]�j�  j�  j  KUubK6j  )��}�(j�  K6j  ]�j�  j�  j  KUubK7j  )��}�(j�  K7j  ]�j�  j�  j  KUubK8j  )��}�(j�  K8j  ]�j�  j�  j  KUubK9j  )��}�(j�  K9j  ]�j�  j�  j  KUubK:j  )��}�(j�  K:j  ]�j�  j�  j  KUubK;j  )��}�(j�  K;j  ]�j�  j�  j  KUubK<j  )��}�(j�  K<j  ]�j�  j�  j  KUubK=j  )��}�(j�  K=j  ]�j�  j�  j  KUubK>j  )��}�(j�  K>j  ]�j�  j�  j  KUubK?j  )��}�(j�  K?j  ]�j�  j�  j  KUubK@j  )��}�(j�  K@j  ]�j�  j�  j  KUubKAj  )��}�(j�  KAj  ]�j�  j�  j  KUubKBj  )��}�(j�  KBj  ]�j�  j�  j  KUubKCj  )��}�(j�  KCj  ]�j�  j�  j  KUubKDj  )��}�(j�  KDj  ]�j�  j�  j  KUubKEj  )��}�(j�  KEj  ]�j�  j�  j  KUubKFj  )��}�(j�  KFj  ]�j�  j�  j  KUubKGj  )��}�(j�  KGj  ]�j�  j�  j  KUubKHj  )��}�(j�  KHj  ]�j�  j�  j  KUubKIj  )��}�(j�  KIj  ]�j�  j�  j  KUubKJj  )��}�(j�  KJj  ]�j�  j�  j  KUubKKj  )��}�(j�  KKj  ]�j�  j�  j  KUubKLj  )��}�(j�  KLj  ]�j�  j�  j  KUubKMj  )��}�(j�  KMj  ]�j�  j�  j  KUubKNj  )��}�(j�  KNj  ]�j�  j�  j  KUubKOj  )��}�(j�  KOj  ]�j�  j�  j  KUubKPj  )��}�(j�  KPj  ]�j�  j�  j  KUubKQj  )��}�(j�  KQj  ]�j�  j�  j  KUubKRj  )��}�(j�  KRj  ]�j�  j�  j  KUubKSj  )��}�(j�  KSj  ]�j�  j�  j  KUubKTj  )��}�(j�  KTj  ]�j�  j�  j  KUubKUj  )��}�(j�  KUj  ]�j�  j�  j  KUubKVj  )��}�(j�  KVj  ]�j�  j�  j  KUubKWj  )��}�(j�  KWj  ]�j�  j�  j  KUubKXj  )��}�(j�  KXj  ]�j�  j�  j  KUubKYj  )��}�(j�  KYj  ]�j�  j�  j  KUubKZj  )��}�(j�  KZj  ]�j�  j�  j  KUubK[j  )��}�(j�  K[j  ]�j�  j�  j  KUubK\j  )��}�(j�  K\j  ]�j�  j�  j  KUubK]j  )��}�(j�  K]j  ]�j�  j�  j  KUubK^j  )��}�(j�  K^j  ]�j�  j�  j  KUubK_j  )��}�(j�  K_j  ]�j�  j�  j  KUubK`j  )��}�(j�  K`j  ]�j�  j�  j  KUubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KUubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KUubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KUubuKV}�(K j  )��}�(j�  K j  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubK	j  )��}�(j�  K	j  ]�j�  j�  j  KVubK
j  )��}�(j�  K
j  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubKj  )��}�(j�  Kj  ]�j�  j�  j  KVubK j  )��}�(j�  K j  ]�j�  j�  j  KVubK!j  )��}�(j�  K!j  ]�j�  j�  j  KVubK"j  )��}�(j�  K"j  ]�j�  j�  j  KVubK#j  )��}�(j�  K#j  ]�j�  j�  j  KVubK$j  )��}�(j�  K$j  ]�j�  j�  j  KVubK%j  )��}�(j�  K%j  ]�j�  j�  j  KVubK&j  )��}�(j�  K&j  ]�j�  j�  j  KVubK'j  )��}�(j�  K'j  ]�j�  j�  j  KVubK(j  )��}�(j�  K(j  ]�j�  j�  j  KVubK)j  )��}�(j�  K)j  ]�j�  j�  j  KVubK*j  )��}�(j�  K*j  ]�j�  j�  j  KVubK+j  )��}�(j�  K+j  ]�j�  j�  j  KVubK,j  )��}�(j�  K,j  ]�j�  j�  j  KVubK-j  )��}�(j�  K-j  ]�j�  j�  j  KVubK.j  )��}�(j�  K.j  ]�j�  j�  j  KVubK/j  )��}�(j�  K/j  ]�j�  j�  j  KVubK0j  )��}�(j�  K0j  ]�j�  j�  j  KVubK1j  )��}�(j�  K1j  ]�j�  j�  j  KVubK2j  )��}�(j�  K2j  ]�j�  j�  j  KVubK3j  )��}�(j�  K3j  ]�j�  j�  j  KVubK4j  )��}�(j�  K4j  ]�j�  j�  j  KVubK5j  )��}�(j�  K5j  ]�j�  j�  j  KVubK6j  )��}�(j�  K6j  ]�j�  j�  j  KVubK7j  )��}�(j�  K7j  ]�j�  j�  j  KVubK8j  )��}�(j�  K8j  ]�j�  j�  j  KVubK9j  )��}�(j�  K9j  ]�j�  j�  j  KVubK:j  )��}�(j�  K:j  ]�j�  j�  j  KVubK;j  )��}�(j�  K;j  ]�j�  j�  j  KVubK<j  )��}�(j�  K<j  ]�j�  j�  j  KVubK=j  )��}�(j�  K=j  ]�j�  j�  j  KVubK>j  )��}�(j�  K>j  ]�j�  j�  j  KVubK?j  )��}�(j�  K?j  ]�j�  j�  j  KVubK@j  )��}�(j�  K@j  ]�j�  j�  j  KVubKAj  )��}�(j�  KAj  ]�j�  j�  j  KVubKBj  )��}�(j�  KBj  ]�j�  j�  j  KVubKCj  )��}�(j�  KCj  ]�j�  j�  j  KVubKDj  )��}�(j�  KDj  ]�j�  j�  j  KVubKEj  )��}�(j�  KEj  ]�j�  j�  j  KVubKFj  )��}�(j�  KFj  ]�j�  j�  j  KVubKGj  )��}�(j�  KGj  ]�j�  j�  j  KVubKHj  )��}�(j�  KHj  ]�j�  j�  j  KVubKIj  )��}�(j�  KIj  ]�j�  j�  j  KVubKJj  )��}�(j�  KJj  ]�j�  j�  j  KVubKKj  )��}�(j�  KKj  ]�j�  j�  j  KVubKLj  )��}�(j�  KLj  ]�j�  j�  j  KVubKMj  )��}�(j�  KMj  ]�j�  j�  j  KVubKNj  )��}�(j�  KNj  ]�j�  j�  j  KVubKOj  )��}�(j�  KOj  ]�j�  j�  j  KVubKPj  )��}�(j�  KPj  ]�j�  j�  j  KVubKQj  )��}�(j�  KQj  ]�j�  j�  j  KVubKRj  )��}�(j�  KRj  ]�j�  j�  j  KVubKSj  )��}�(j�  KSj  ]�j�  j�  j  KVubKTj  )��}�(j�  KTj  ]�j�  j�  j  KVubKUj  )��}�(j�  KUj  ]�j�  j�  j  KVubKVj  )��}�(j�  KVj  ]�j�  j�  j  KVubKWj  )��}�(j�  KWj  ]�j�  j�  j  KVubKXj  )��}�(j�  KXj  ]�j�  j�  j  KVubKYj  )��}�(j�  KYj  ]�j�  j�  j  KVubKZj  )��}�(j�  KZj  ]�j�  j�  j  KVubK[j  )��}�(j�  K[j  ]�j�  j�  j  KVubK\j  )��}�(j�  K\j  ]�j�  j�  j  KVubK]j  )��}�(j�  K]j  ]�j�  j�  j  KVubK^j  )��}�(j�  K^j  ]�j�  j�  j  KVubK_j  )��}�(j�  K_j  ]�j�  j�  j  KVubK`j  )��}�(j�  K`j  ]�j�  j�  j  KVubKaj  )��}�(�       j�  Kaj  ]�j�  j�  j  KVubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KVubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KVubuKW}�(K j  )��}�(j�  K j  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubK	j  )��}�(j�  K	j  ]�j�  j�  j  KWubK
j  )��}�(j�  K
j  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubKj  )��}�(j�  Kj  ]�j�  j�  j  KWubK j  )��}�(j�  K j  ]�j�  j�  j  KWubK!j  )��}�(j�  K!j  ]�j�  j�  j  KWubK"j  )��}�(j�  K"j  ]�j�  j�  j  KWubK#j  )��}�(j�  K#j  ]�j�  j�  j  KWubK$j  )��}�(j�  K$j  ]�j�  j�  j  KWubK%j  )��}�(j�  K%j  ]�j�  j�  j  KWubK&j  )��}�(j�  K&j  ]�j�  j�  j  KWubK'j  )��}�(j�  K'j  ]�j�  j�  j  KWubK(j  )��}�(j�  K(j  ]�j�  j�  j  KWubK)j  )��}�(j�  K)j  ]�j�  j�  j  KWubK*j  )��}�(j�  K*j  ]�j�  j�  j  KWubK+j  )��}�(j�  K+j  ]�j�  j�  j  KWubK,j  )��}�(j�  K,j  ]�j�  j�  j  KWubK-j  )��}�(j�  K-j  ]�j�  j�  j  KWubK.j  )��}�(j�  K.j  ]�j�  j�  j  KWubK/j  )��}�(j�  K/j  ]�j�  j�  j  KWubK0j  )��}�(j�  K0j  ]�j�  j�  j  KWubK1j  )��}�(j�  K1j  ]�j�  j�  j  KWubK2j  )��}�(j�  K2j  ]�j�  j�  j  KWubK3j  )��}�(j�  K3j  ]�j�  j�  j  KWubK4j  )��}�(j�  K4j  ]�j�  j�  j  KWubK5j  )��}�(j�  K5j  ]�j�  j�  j  KWubK6j  )��}�(j�  K6j  ]�j�  j�  j  KWubK7j  )��}�(j�  K7j  ]�j�  j�  j  KWubK8j  )��}�(j�  K8j  ]�j�  j�  j  KWubK9j  )��}�(j�  K9j  ]�j�  j�  j  KWubK:j  )��}�(j�  K:j  ]�j�  j�  j  KWubK;j  )��}�(j�  K;j  ]�j�  j�  j  KWubK<j  )��}�(j�  K<j  ]�j�  j�  j  KWubK=j  )��}�(j�  K=j  ]�j�  j�  j  KWubK>j  )��}�(j�  K>j  ]�j�  j�  j  KWubK?j  )��}�(j�  K?j  ]�j�  j�  j  KWubK@j  )��}�(j�  K@j  ]�j�  j�  j  KWubKAj  )��}�(j�  KAj  ]�j�  j�  j  KWubKBj  )��}�(j�  KBj  ]�j�  j�  j  KWubKCj  )��}�(j�  KCj  ]�j�  j�  j  KWubKDj  )��}�(j�  KDj  ]�j�  j�  j  KWubKEj  )��}�(j�  KEj  ]�j�  j�  j  KWubKFj  )��}�(j�  KFj  ]�j�  j�  j  KWubKGj  )��}�(j�  KGj  ]�j�  j�  j  KWubKHj  )��}�(j�  KHj  ]�j�  j�  j  KWubKIj  )��}�(j�  KIj  ]�j�  j�  j  KWubKJj  )��}�(j�  KJj  ]�j�  j�  j  KWubKKj  )��}�(j�  KKj  ]�j�  j�  j  KWubKLj  )��}�(j�  KLj  ]�j�  j�  j  KWubKMj  )��}�(j�  KMj  ]�j�  j�  j  KWubKNj  )��}�(j�  KNj  ]�j�  j�  j  KWubKOj  )��}�(j�  KOj  ]�j�  j�  j  KWubKPj  )��}�(j�  KPj  ]�j�  j�  j  KWubKQj  )��}�(j�  KQj  ]�j�  j�  j  KWubKRj  )��}�(j�  KRj  ]�j�  j�  j  KWubKSj  )��}�(j�  KSj  ]�j�  j�  j  KWubKTj  )��}�(j�  KTj  ]�j�  j�  j  KWubKUj  )��}�(j�  KUj  ]�j�  j�  j  KWubKVj  )��}�(j�  KVj  ]�j�  j�  j  KWubKWj  )��}�(j�  KWj  ]�j�  j�  j  KWubKXj  )��}�(j�  KXj  ]�j�  j�  j  KWubKYj  )��}�(j�  KYj  ]�j�  j�  j  KWubKZj  )��}�(j�  KZj  ]�j�  j�  j  KWubK[j  )��}�(j�  K[j  ]�j�  j�  j  KWubK\j  )��}�(j�  K\j  ]�j�  j�  j  KWubK]j  )��}�(j�  K]j  ]�j�  j�  j  KWubK^j  )��}�(j�  K^j  ]�j�  j�  j  KWubK_j  )��}�(j�  K_j  ]�j�  j�  j  KWubK`j  )��}�(j�  K`j  ]�j�  j�  j  KWubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KWubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KWubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KWubuKX}�(K j  )��}�(j�  K j  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubK	j  )��}�(j�  K	j  ]�j�  j�  j  KXubK
j  )��}�(j�  K
j  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubKj  )��}�(j�  Kj  ]�j�  j�  j  KXubK j  )��}�(j�  K j  ]�j�  j�  j  KXubK!j  )��}�(j�  K!j  ]�j�  j�  j  KXubK"j  )��}�(j�  K"j  ]�j�  j�  j  KXubK#j  )��}�(j�  K#j  ]�j�  j�  j  KXubK$j  )��}�(j�  K$j  ]�j�  j�  j  KXubK%j  )��}�(j�  K%j  ]�j�  j�  j  KXubK&j  )��}�(j�  K&j  ]�j�  j�  j  KXubK'j  )��}�(j�  K'j  ]�j�  j�  j  KXubK(j  )��}�(j�  K(j  ]�j�  j�  j  KXubK)j  )��}�(j�  K)j  ]�j�  j�  j  KXubK*j  )��}�(j�  K*j  ]�j�  j�  j  KXubK+j  )��}�(j�  K+j  ]�j�  j�  j  KXubK,j  )��}�(j�  K,j  ]�j�  j�  j  KXubK-j  )��}�(j�  K-j  ]�j�  j�  j  KXubK.j  )��}�(j�  K.j  ]�j�  j�  j  KXubK/j  )��}�(j�  K/j  ]�j�  j�  j  KXubK0j  )��}�(j�  K0j  ]�j�  j�  j  KXubK1j  )��}�(j�  K1j  ]�j�  j�  j  KXubK2j  )��}�(j�  K2j  ]�j�  j�  j  KXubK3j  )��}�(j�  K3j  ]�j�  j�  j  KXubK4j  )��}�(j�  K4j  ]�j�  j�  j  KXubK5j  )��}�(j�  K5j  ]�j�  j�  j  KXubK6j  )��}�(j�  K6j  ]�j�  j�  j  KXubK7j  )��}�(j�  K7j  ]�j�  j�  j  KXubK8j  )��}�(j�  K8j  ]�j�  j�  j  KXubK9j  )��}�(j�  K9j  ]�j�  j�  j  KXubK:j  )��}�(j�  K:j  ]�j�  j�  j  KXubK;j  )��}�(j�  K;j  ]�j�  j�  j  KXubK<j  )��}�(j�  K<j  ]�j�  j�  j  KXubK=j  )��}�(j�  K=j  ]�j�  j�  j  KXubK>j  )��}�(j�  K>j  ]�j�  j�  j  KXubK?j  )��}�(j�  K?j  ]�j�  j�  j  KXubK@j  )��}�(j�  K@j  ]�j�  j�  j  KXubKAj  )��}�(j�  KAj  ]�j�  j�  j  KXubKBj  )��}�(j�  KBj  ]�j�  j�  j  KXubKCj  )��}�(j�  KCj  ]�j�  j�  j  KXubKDj  )��}�(j�  KDj  ]�j�  j�  j  KXubKEj  )��}�(j�  KEj  ]�j�  j�  j  KXubKFj  )��}�(j�  KFj  ]�j�  j�  j  KXubKGj  )��}�(j�  KGj  ]�j�  j�  j  KXubKHj  )��}�(j�  KHj  ]�j�  j�  j  KXubKIj  )��}�(j�  KIj  ]�j�  j�  j  KXubKJj  )��}�(j�  KJj  ]�j�  j�  j  KXubKKj  )��}�(j�  KKj  ]�j�  j�  j  KXubKLj  )��}�(j�  KLj  ]�j�  j�  j  KXubKMj  )��}�(j�  KMj  ]�j�  j�  j  KXubKNj  )��}�(j�  KNj  ]�j�  j�  j  KXubKOj  )��}�(j�  KOj  ]�j�  j�  j  KXubKPj  )��}�(j�  KPj  ]�j�  j�  j  KXubKQj  )��}�(j�  KQj  ]�j�  j�  j  KXubKRj  )��}�(j�  KRj  ]�j�  j�  j  KXubKSj  )��}�(j�  KSj  ]�j�  j�  j  KXubKTj  )��}�(j�  KTj  ]�j�  j�  j  KXubKUj  )��}�(j�  KUj  ]�j�  j�  j  KXubKVj  )��}�(j�  KVj  ]�j�  j�  j  KXubKWj  )��}�(j�  KWj  ]�j�  j�  j  KXubKXj  )��}�(j�  KXj  ]�j�  j�  j  KXubKYj  )��}�(j�  KYj  ]�j�  j�  j  KXubKZj  )��}�(j�  KZj  ]�j�  j�  j  KXubK[j  )��}�(j�  K[j  ]�j�  j�  j  KXubK\j  )��}�(j�  K\j  ]�j�  j�  j  KXubK]j  )��}�(j�  K]j  ]�j�  j�  j  KXubK^j  )��}�(j�  K^j  ]�j�  j�  j  KXubK_j  )��}�(j�  K_j  ]�j�  j�  j  KXubK`j  )��}�(j�  K`j  ]�j�  j�  j  KXubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KXubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KXubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KXubuKY}�(K j  )��}�(j�  K j  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubK	j  )��}�(j�  K	j  ]�j�  j�  j  KYubK
j  )��}�(j�  K
j  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubKj  )��}�(j�  Kj  ]�j�  j�  j  KYubK j  )��}�(j�  K j  ]�j�  j�  j  KYubK!j  )��}�(j�  K!j  ]�j�  j�  j  KYubK"j  )��}�(j�  K"j  ]�j�  j�  j  KYubK#j  )��}�(j�  K#j  ]�j�  j�  j  KYubK$j  )��}�(j�  K$j  ]�j�  j�  j  KYubK%j  )��}�(j�  K%j  ]�j�  j�  j  KYubK&j  )��}�(j�  K&j  ]�j�  j�  j  KYubK'j  )��}�(j�  K'j  ]�j�  j�  j  KYubK(j  )��}�(j�  K(j  ]�j�  j�  j  KYubK)j  )��}�(j�  K)j  ]�j�  j�  j  KYubK*j  )��}�(j�  K*j  ]�j�  j�  j  KYubK+j  )��}�(j�  K+j  ]�j�  j�  j  KYubK,j  )��}�(j�  K,j  ]�j�  j�  j  KYubK-j  )��}�(j�  K-j  ]�j�  j�  j  KYubK.j  )��}�(j�  K.j  ]�j�  j�  j  KYubK/j  )��}�(j�  K/j  ]�j�  j�  j  KYubK0j  )��}�(j�  K0j  ]�j�  j�  j  KYubK1j  )��}�(j�  K1j  ]�j�  j�  j  KYubK2j  )��}�(j�  K2j  ]�j�  j�  j  KYubK3j  )��}�(j�  K3j  ]�j�  j�  j  KYubK4j  )��}�(j�  K4j  ]�j�  j�  j  KYubK5j  )��}�(j�  K5j  ]�j�  j�  j  KYubK6j  )��}�(j�  K6j  ]�j�  j�  j  KYubK7j  )��}�(j�  K7j  ]�j�  j�  j  KYubK8j  )��}�(j�  K8j  ]�j�  j�  j  KYubK9j  )��}�(j�  K9j  ]�j�  j�  j  KYubK:j  )��}�(j�  K:j  ]�j�  j�  j  KYubK;j  )��}�(j�  K;j  ]�j�  j�  j  KYubK<j  )��}�(j�  K<j  ]�j�  j�  j  KYubK=j  )��}�(j�  K=j  ]�j�  j�  j  KYubK>j  )��}�(j�  K>j  ]�j�  j�  j  KYubK?j  )��}�(j�  K?j  ]�j�  j�  j  KYubK@j  )��}�(j�  K@j  ]�j�  j�  j  KYubKAj  )��}�(j�  KAj  ]�j�  j�  j  KYubKBj  )��}�(j�  KBj  ]�j�  j�  j  KYubKCj  )��}�(j�  KCj  ]�j�  j�  j  KYubKDj  )��}�(j�  KDj  ]�j�  j�  j  KYubKEj  )��}�(j�  KEj  ]�j�  j�  j  KYubKFj  )��}�(j�  KFj  ]�j�  j�  j  KYubKGj  )��}�(j�  KGj  ]�j�  j�  j  KYubKHj  )��}�(j�  KHj  ]�j�  j�  j  KYubKIj  )��}�(j�  KIj  ]�j�  j�  j  KYubKJj  )��}�(j�  KJj  ]�j�  j�  j  KYubKKj  )��}�(j�  KKj  ]�j�  j�  j  KYubKLj  )��}�(j�  KLj  ]�j�  j�  j  KYubKMj  )��}�(j�  KMj  ]�j�  j�  j  KYubKNj  )��}�(j�  KNj  ]�j�  j�  j  KYubKOj  )��}�(j�  KOj  ]�j�  j�  j  KYubKPj  )��}�(j�  KPj  ]�j�  j�  j  KYubKQj  )��}�(j�  KQj  ]�j�  j�  j  KYubKRj  )��}�(j�  KRj  ]�j�  j�  j  KYubKSj  )��}�(j�  KSj  ]�j�  j�  j  KYubKTj  )��}�(j�  KTj  ]�j�  j�  j  KYubKUj  )��}�(j�  KUj  ]�j�  j�  j  KYubKVj  )��}�(j�  KVj  ]�j�  j�  j  KYubKWj  )��}�(j�  KWj  ]�j�  j�  j  KYubKXj  )��}�(j�  KXj  ]�j�  j�  j  KYubKYj  )��}�(j�  KYj  ]�j�  j�  j  KYubKZj  )��}�(j�  KZj  ]�j�  j�  j  KYubK[j  )��}�(j�  K[j  ]�j�  j�  j  KYubK\j  )��}�(j�  K\j  ]�j�  j�  j  KYubK]j  )��}�(j�  K]j  ]�j�  j�  j  KYubK^j  )��}�(j�  K^j  ]�j�  j�  j  KYubK_j  )��}�(j�  K_j  ]�j�  j�  j  KYubK`j  )��}�(j�  K`j  ]�j�  j�  j  KYubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KYubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KYubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KYubuKZ}�(K j  )��}�(j�  K j  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubK	j  )��}�(j�  K	j  ]�j�  j�  j  KZubK
j  )��}�(j�  K
j  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubKj  )��}�(j�  Kj  ]�j�  j�  j  KZubK j  )��}�(j�  K j  ]�j�  j�  j  KZubK!j  )��}�(j�  K!j  ]�j�  j�  j  KZubK"j  )��}�(j�  K"j  ]�j�  j�  j  KZubK#j  )��}�(j�  K#j  ]�j�  j�  j  KZubK$j  )��}�(j�  K$j  ]�j�  j�  j  KZubK%j  )��}�(j�  K%j  ]�j�  j�  j  KZubK&j  )��}�(j�  K&j  ]�j�  j�  j  KZubK'j  )��}�(j�  K'j  ]�j�  j�  j  KZubK(j  )��}�(j�  K(j  ]�j�  j�  j  KZubK)j  )��}�(j�  K)j  ]�j�  j�  j  KZubK*j  )��}�(j�  K*j  ]�j�  j�  j  KZubK+j  )��}�(j�  K+j  ]�j�  j�  j  KZubK,j  )��}�(j�  K,j  ]�j�  j�  j  KZubK-j  )��}�(j�  K-j  ]�j�  j�  j  KZubK.j  )��}�(j�  K.j  ]�j�  j�  j  KZubK/j  )��}�(j�  K/j  ]�j�  j�  j  KZubK0j  )��}�(j�  K0j  ]�j�  j�  j  KZubK1j  )��}�(j�  K1j  ]�j�  j�  j  KZubK2j  )��}�(j�  K2j  ]�j�  j�  j  KZubK3j  )��}�(j�  K3j  ]�j�  j�  j  KZubK4j  )��}�(j�  K4j  ]�j�  j�  j  KZubK5j  )��}�(j�  K5j  ]�j�  j�  j  KZubK6j  )��}�(j�  K6j  ]�j�  j�  j  KZubK7j  )��}�(j�  K7j  ]�j�  j�  j  KZubK8j  )��}�(j�  K8j  ]�j�  j�  j  KZubK9j  )��}�(j�  K9j  ]�j�  j�  j  KZubK:j  )��}�(j�  K:j  ]�j�  j�  j  KZubK;j  )��}�(j�  K;j  ]�j�  j�  j  KZubK<j  )��}�(j�  K<j  ]�j�  j�  j  KZubK=j  )��}�(j�  K=j  ]�j�  j�  j  KZubK>j  )��}�(j�  K>j  ]�j�  j�  j  KZubK?j  )��}�(j�  K?j  ]�j�  j�  j  KZubK@j  )��}�(j�  K@j  ]�j�  j�  j  KZubKAj  )��}�(j�  KAj  ]�j�  j�  j  KZubKBj  )��}�(j�  KBj  ]�j�  j�  j  KZubKCj  )��}�(j�  KCj  ]�j�  j�  j  KZubKDj  )��}�(j�  KDj  ]�j�  j�  j  KZubKEj  )��}�(j�  KEj  ]�j�  j�  j  KZubKFj  )��}�(j�  KFj  ]�j�  j�  j  KZubKGj  )��}�(j�  KGj  ]�j�  j�  j  KZubKHj  )��}�(j�  KHj  ]�j�  j�  j  KZubKIj  )��}�(j�  KIj  ]�j�  j�  j  KZubKJj  )��}�(j�  KJj  ]�j�  j�  j  KZubKKj  )��}�(j�  KKj  ]�j�  j�  j  KZubKLj  )��}�(j�  KLj  ]�j�  j�  j  KZubKMj  )��}�(j�  KMj  ]�j�  j�  j  KZubKNj  )��}�(j�  KNj  ]�j�  j�  j  KZubKOj  )��}�(j�  KOj  ]�j�  j�  j  KZubKPj  )��}�(j�  KPj  ]�j�  j�  j  KZubKQj  )��}�(j�  KQj  ]�j�  j�  j  KZubKRj  )��}�(j�  KRj  ]�j�  j�  j  KZubKSj  )��}�(j�  KSj  ]�j�  j�  j  KZubKTj  )��}�(j�  KTj  ]�j�  j�  j  KZubKUj  )��}�(j�  KUj  ]�j�  j�  j  KZubKVj  )��}�(j�  KVj  ]�j�  j�  j  KZubKWj  )��}�(j�  KWj  ]�j�  j�  j  KZubKXj  )��}�(j�  KXj  ]�j�  j�  j  KZubKYj  )��}�(j�  KYj  ]�j�  j�  j  KZubKZj  )��}�(j�  KZj  ]�j�  j�  j  KZubK[j  )��}�(j�  K[j  ]�j�  j�  j  KZubK\j  )��}�(j�  K\j  ]�j�  j�  j  KZubK]j  )��}�(j�  K]j  ]�j�  j�  j  KZubK^j  )��}�(j�  K^j  ]�j�  j�  j  KZubK_j  )��}�(j�  K_j  ]�j�  j�  j  KZubK`j  )��}�(j�  K`j  ]�j�  j�  j  KZubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KZubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KZubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KZubuK[}�(K j  )��}�(j�  K j  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K[ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubKj  )��}�(j�  Kj  ]�j�  j�  j  K[ubK j  )��}�(j�  K j  ]�j�  j�  j  K[ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K[ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K[ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K[ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K[ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K[ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K[ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K[ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K[ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K[ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K[ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K[ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K[ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K[ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K[ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K[ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K[ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K[ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K[ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K[ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K[ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K[ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K[ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K[ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K[ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K[ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K[ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K[ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K[ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K[ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K[ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K[ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K[ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K[ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K[ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K[ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K[ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K[ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K[ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K[ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K[ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K[ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K[ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K[ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K[ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K[ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K[ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K[ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K[ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K[ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K[ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K[ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K[ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K[ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K[ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K[ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K[ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K[ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K[ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K[ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K[ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K[ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K[ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K[ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K[ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K[ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K[ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K[ubuK\}�(K j  )��}�(j�  K j  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K\ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubKj  )��}�(j�  Kj  ]�j�  j�  j  K\ubK j  )��}�(j�  K j  ]�j�  j�  j  K\ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K\ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K\ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K\ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K\ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K\ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K\ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K\ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K\ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K\ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K\ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K\ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K\ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K\ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K\ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K\ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K\ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K\ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K\ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K\ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K\ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K\ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K\ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K\ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K\ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K\ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K\ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K\ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K\ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K\ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K\ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K\ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K\ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K\ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K\ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K\ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K\ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K\ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K\ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K\ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K\ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K\ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K\ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K\ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K\ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K\ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K\ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K\ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K\ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K\ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K\ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K\ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K\ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K\ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K\ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K\ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K\ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K\ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K\ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K\ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K\ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K\ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K\ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K\ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K\ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K\ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K\ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K\ubuK]}�(K j  )��}�(j�  K j  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K]ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubKj  )��}�(j�  Kj  ]�j�  j�  j  K]ubK j  )��}�(j�  K j  ]�j�  j�  j  K]ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K]ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K]ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K]ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K]ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K]ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K]ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K]ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K]ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K]ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K]ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K]ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K]ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K]ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K]ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K]ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K]ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K]ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K]ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K]ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K]ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K]ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K]ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K]ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K]ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K]ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K]ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K]ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K]ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K]ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K]ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K]ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K]ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K]ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K]ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K]ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K]ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K]ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K]ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K]ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K]ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K]ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K]ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K]ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K]ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K]ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K]ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K]ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K]ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K]ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K]ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K]ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K]ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K]ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K]ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K]ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K]ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K]ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K]ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K]ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K]ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K]ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K]ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K]ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K]ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K]ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K]ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K]ubuK^}�(K j  )��}�(j�  K j  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K^ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubKj  )��}�(j�  Kj  ]�j�  j�  j  K^ubK j  )��}�(j�  K j  ]�j�  j�  j  K^ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K^ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K^ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K^ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K^ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K^ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K^ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K^ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K^ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K^ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K^ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K^ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K^ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K^ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K^ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K^ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K^ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K^ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K^ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K^ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K^ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K^ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K^ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K^ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K^ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K^ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K^ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K^ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K^ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K^ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K^ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K^ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K^ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K^ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K^ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K^ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K^ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K^ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K^ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K^ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K^ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K^ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K^ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K^ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K^ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K^ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K^ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K^ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K^ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K^ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K^ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K^ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K^ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K^ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K^ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K^ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K^ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K^ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K^ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K^ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K^ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K^ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K^ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K^ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K^ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K^ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K^ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K^ubuK_}�(K j  )��}�(j�  K j  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K_ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubKj  )��}�(j�  Kj  ]�j�  j�  j  K_ubK j  )��}�(j�  K j  ]�j�  j�  j  K_ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K_ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K_ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K_ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K_ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K_ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K_ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K_ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K_ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K_ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K_ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K_ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K_ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K_ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K_ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K_ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K_ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K_ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K_ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K_ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K_ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K_ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K_ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K_ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K_ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K_ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K_ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K_ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K_ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K_ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K_ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K_ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K_ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K_ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K_ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K_ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K_ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K_ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K_ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K_ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K_ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K_ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K_ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K_ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K_ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K_ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K_ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K_ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K_ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K_ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K_ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K_ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K_ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K_ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K_ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K_ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K_ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K_ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K_ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K_ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K_ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K_ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K_ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K_ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K_ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K_ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K_ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K_ubuK`}�(K j  )��}�(j�  K j  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubK	j  )��}�(j�  K	j  ]�j�  j�  j  K`ubK
j  )��}�(j�  K
j  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubKj  )��}�(j�  Kj  ]�j�  j�  j  K`ubK j  )��}�(j�  K j  ]�j�  j�  j  K`ubK!j  )��}�(j�  K!j  ]�j�  j�  j  K`ubK"j  )��}�(j�  K"j  ]�j�  j�  j  K`ubK#j  )��}�(j�  K#j  ]�j�  j�  j  K`ubK$j  )��}�(j�  K$j  ]�j�  j�  j  K`ubK%j  )��}�(j�  K%j  ]�j�  j�  j  K`ubK&j  )��}�(j�  K&j  ]�j�  j�  j  K`ubK'j  )��}�(j�  K'j  ]�j�  j�  j  K`ubK(j  )��}�(j�  K(j  ]�j�  j�  j  K`ubK)j  )��}�(j�  K)j  ]�j�  j�  j  K`ubK*j  )��}�(j�  K*j  ]�j�  j�  j  K`ubK+j  )��}�(j�  K+j  ]�j�  j�  j  K`ubK,j  )��}�(j�  K,j  ]�j�  j�  j  K`ubK-j  )��}�(j�  K-j  ]�j�  j�  j  K`ubK.j  )��}�(j�  K.j  ]�j�  j�  j  K`ubK/j  )��}�(j�  K/j  ]�j�  j�  j  K`ubK0j  )��}�(j�  K0j  ]�j�  j�  j  K`ubK1j  )��}�(j�  K1j  ]�j�  j�  j  K`ubK2j  )��}�(j�  K2j  ]�j�  j�  j  K`ubK3j  )��}�(j�  K3j  ]�j�  j�  j  K`ubK4j  )��}�(j�  K4j  ]�j�  j�  j  K`ubK5j  )��}�(j�  K5j  ]�j�  j�  j  K`ubK6j  )��}�(j�  K6j  ]�j�  j�  j  K`ubK7j  )��}�(j�  K7j  ]�j�  j�  j  K`ubK8j  )��}�(j�  K8j  ]�j�  j�  j  K`ubK9j  )��}�(j�  K9j  ]�j�  j�  j  K`ubK:j  )��}�(j�  K:j  ]�j�  j�  j  K`ubK;j  )��}�(j�  K;j  ]�j�  j�  j  K`ubK<j  )��}�(j�  K<j  ]�j�  j�  j  K`ubK=j  )��}�(j�  K=j  ]�j�  j�  j  K`ubK>j  )��}�(j�  K>j  ]�j�  j�  j  K`ubK?j  )��}�(j�  K?j  ]�j�  j�  j  K`ubK@j  )��}�(j�  K@j  ]�j�  j�  j  K`ubKAj  )��}�(j�  KAj  ]�j�  j�  j  K`ubKBj  )��}�(j�  KBj  ]�j�  j�  j  K`ubKCj  )��}�(j�  KCj  ]�j�  j�  j  K`ubKDj  )��}�(j�  KDj  ]�j�  j�  j  K`ubKEj  )��}�(j�  KEj  ]�j�  j�  j  K`ubKFj  )��}�(j�  KFj  ]�j�  j�  j  K`ubKGj  )��}�(j�  KGj  ]�j�  j�  j  K`ubKHj  )��}�(j�  KHj  ]�j�  j�  j  K`ubKIj  )��}�(j�  KIj  ]�j�  j�  j  K`ubKJj  )��}�(j�  KJj  ]�j�  j�  j  K`ubKKj  )��}�(j�  KKj  ]�j�  j�  j  K`ubKLj  )��}�(j�  KLj  ]�j�  j�  j  K`ubKMj  )��}�(j�  KMj  ]�j�  j�  j  K`ubKNj  )��}�(j�  KNj  ]�j�  j�  j  K`ubKOj  )��}�(j�  KOj  ]�j�  j�  j  K`ubKPj  )��}�(j�  KPj  ]�j�  j�  j  K`ubKQj  )��}�(j�  KQj  ]�j�  j�  j  K`ubKRj  )��}�(j�  KRj  ]�j�  j�  j  K`ubKSj  )��}�(j�  KSj  ]�j�  j�  j  K`ubKTj  )��}�(j�  KTj  ]�j�  j�  j  K`ubKUj  )��}�(j�  KUj  ]�j�  j�  j  K`ubKVj  )��}�(j�  KVj  ]�j�  j�  j  K`ubKWj  )��}�(j�  KWj  ]�j�  j�  j  K`ubKXj  )��}�(j�  KXj  ]�j�  j�  j  K`ubKYj  )��}�(j�  KYj  ]�j�  j�  j  K`ubKZj  )��}�(j�  KZj  ]�j�  j�  j  K`ubK[j  )��}�(j�  K[j  ]�j�  j�  j  K`ubK\j  )��}�(j�  K\j  ]�j�  j�  j  K`ubK]j  )��}�(j�  K]j  ]�j�  j�  j  K`ubK^j  )��}�(j�  K^j  ]�j�  j�  j  K`ubK_j  )��}�(j�  K_j  ]�j�  j�  j  K`ubK`j  )��}�(j�  K`j  ]�j�  j�  j  K`ubKaj  )��}�(j�  Kaj  ]�j�  j�  j  K`ubKbj  )��}�(j�  Kbj  ]�j�  j�  j  K`ubKcj  )��}�(j�  Kcj  ]�j�  j�  j  K`ubuKa}�(K j  )��}�(j�  K j  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubK	j  )��}�(j�  K	j  ]�j�  j�  j  KaubK
j  )��}�(j�  K
j  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubKj  )��}�(j�  Kj  ]�j�  j�  j  KaubK j  )��}�(j�  K j  ]�j�  j�  j  KaubK!j  )��}�(j�  K!j  ]�j�  j�  j  KaubK"j  )��}�(j�  K"j  ]�j�  j�  j  KaubK#j  )��}�(j�  K#j  ]�j�  j�  j  KaubK$j  )��}�(j�  K$j  ]�j�  j�  j  KaubK%j  )��}�(j�  K%j  ]�j�  j�  j  KaubK&j  )��}�(j�  K&j  ]�j�  j�  j  KaubK'j  )��}�(j�  K'j  ]�j�  j�  j  KaubK(j  )��}�(j�  K(j  ]�j�  j�  j  KaubK)j  )��}�(j�  K)j  ]�j�  j�  j  KaubK*j  )��}�(j�  K*j  ]�j�  j�  j  KaubK+j  )��}�(j�  K+j  ]�j�  j�  j  KaubK,j  )��}�(j�  K,j  ]�j�  j�  j  KaubK-j  )��}�(j�  K-j  ]�j�  j�  j  KaubK.j  )��}�(j�  K.j  ]�j�  j�  j  KaubK/j  )��}�(j�  K/j  ]�j�  j�  j  KaubK0j  )��}�(j�  K0j  ]�j�  j�  j  KaubK1j  )��}�(j�  K1j  ]�j�  j�  j  KaubK2j  )��}�(j�  K2j  ]�j�  j�  j  KaubK3j  )��}�(j�  K3j  ]�j�  j�  j  KaubK4j  )��}�(j�  K4j  ]�j�  j�  j  KaubK5j  )��}�(j�  K5j  ]�j�  j�  j  KaubK6j  )��}�(j�  K6j  ]�j�  j�  j  KaubK7j  )��}�(j�  K7j  ]�j�  j�  j  KaubK8j  )��}�(j�  K8j  ]�j�  j�  j  KaubK9j  )��}�(j�  K9j  ]�j�  j�  j  KaubK:j  )��}�(j�  K:j  ]�j�  j�  j  KaubK;j  )��}�(j�  K;j  ]�j�  j�  j  KaubK<j  )��}�(j�  K<j  ]�j�  j�  j  KaubK=j  )��}�(j�  K=j  ]�j�  j�  j  KaubK>j  )��}�(j�  K>j  ]�j�  j�  j  KaubK?j  )��}�(j�  K?j  ]�j�  j�  j  KaubK@j  )��}�(j�  K@j  ]�j�  j�  j  KaubKAj  )��}�(j�  KAj  ]�j�  j�  j  KaubKBj  )��}�(j�  KBj  ]�j�  j�  j  KaubKCj  )��}�(j�  KCj  ]�j�  j�  j  KaubKDj  )��}�(j�  KDj  ]�j�  j�  j  KaubKEj  )��}�(j�  KEj  ]�j�  j�  j  KaubKFj  )��}�(j�  KFj  ]�j�  j�  j  KaubKGj  )��}�(j�  KGj  ]�j�  j�  j  KaubKHj  )��}�(j�  KHj  ]�j�  j�  j  KaubKIj  )��}�(j�  KIj  ]�j�  j�  j  KaubKJj  )��}�(j�  KJj  ]�j�  j�  j  KaubKKj  )��}�(j�  KKj  ]�j�  j�  j  KaubKLj  )��}�(j�  KLj  ]�j�  j�  j  KaubKMj  )��}�(j�  KMj  ]�j�  j�  j  KaubKNj  )��}�(j�  KNj  ]�j�  j�  j  KaubKOj  )��}�(j�  KOj  ]�j�  j�  j  KaubKPj  )��}�(j�  KPj  ]�j�  j�  j  KaubKQj  )��}�(j�  KQj  ]�j�  j�  j  KaubKRj  )��}�(j�  KRj  ]�j�  j�  j  KaubKSj  )��}�(j�  KSj  ]�j�  j�  j  KaubKTj  )��}�(j�  KTj  ]�j�  j�  j  KaubKUj  )��}�(j�  KUj  ]�j�  j�  j  KaubKVj  )��}�(j�  KVj  ]�j�  j�  j  KaubKWj  )��}�(j�  KWj  ]�j�  j�  j  KaubKXj  )��}�(j�  KXj  ]�j�  j�  j  KaubKYj  )��}�(j�  KYj  ]�j�  j�  j  KaubKZj  )��}�(j�  KZj  ]�j�  j�  j  KaubK[j  )��}�(j�  K[j  ]�j�  j�  j  KaubK\j  )��}�(j�  K\j  ]�j�  j�  j  KaubK]j  )��}�(j�  K]j  ]�j�  j�  j  KaubK^j  )��}�(j�  K^j  ]�j�  j�  j  KaubK_j  )��}�(j�  K_j  ]�j�  j�  j  KaubK`j  )��}�(j�  K`j  ]�j�  j�  j  KaubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KaubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KaubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KaubuKb}�(K j  )��}�(j�  K j  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubK	j  )��}�(j�  K	j  ]�j�  j�  j  KbubK
j  )��}�(j�  K
j  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubKj  )��}�(j�  Kj  ]�j�  j�  j  KbubK j  )��}�(j�  K j  ]�j�  j�  j  KbubK!j  )��}�(j�  K!j  ]�j�  j�  j  KbubK"j  )��}�(j�  K"j  ]�j�  j�  j  KbubK#j  )��}�(j�  K#j  ]�j�  j�  j  KbubK$j  )��}�(j�  K$j  ]�j�  j�  j  KbubK%j  )��}�(j�  K%j  ]�j�  j�  j  KbubK&j  )��}�(j�  K&j  ]�j�  j�  j  KbubK'j  )��}�(j�  K'j  ]�j�  j�  j  KbubK(j  )��}�(j�  K(j  ]�j�  j�  j  KbubK)j  )��}�(j�  K)j  ]�j�  j�  j  KbubK*j  )��}�(j�  K*j  ]�j�  j�  j  KbubK+j  )��}�(j�  K+j  ]�j�  j�  j  KbubK,j  )��}�(j�  K,j  ]�j�  j�  j  KbubK-j  )��}�(j�  K-j  ]�j�  j�  j  KbubK.j  )��}�(j�  K.j  ]�j�  j�  j  KbubK/j  )��}�(j�  K/j  ]�j�  j�  j  KbubK0j  )��}�(j�  K0j  ]�j�  j�  j  KbubK1j  )��}�(j�  K1j  ]�j�  j�  j  KbubK2j  )��}�(j�  K2j  ]�j�  j�  j  KbubK3j  )��}�(j�  K3j  ]�j�  j�  j  KbubK4j  )��}�(j�  K4j  ]�j�  j�  j  KbubK5j  )��}�(j�  K5j  ]�j�  j�  j  KbubK6j  )��}�(j�  K6j  ]�j�  j�  j  KbubK7j  )��}�(j�  K7j  ]�j�  j�  j  KbubK8j  )��}�(j�  K8j  ]�j�  j�  j  KbubK9j  )��}�(j�  K9j  ]�j�  j�  j  KbubK:j  )��}�(j�  K:j  ]�j�  j�  j  KbubK;j  )��}�(j�  K;j  ]�j�  j�  j  KbubK<j  )��}�(j�  K<j  ]�j�  j�  j  KbubK=j  )��}�(j�  K=j  ]�j�  j�  j  KbubK>j  )��}�(j�  K>j  ]�j�  j�  j  KbubK?j  )��}�(j�  K?j  ]�j�  j�  j  KbubK@j  )��}�(j�  K@j  ]�j�  j�  j  KbubKAj  )��}�(j�  KAj  ]�j�  j�  j  KbubKBj  )��}�(j�  KBj  ]�j�  j�  j  KbubKCj  )��}�(j�  KCj  ]�j�  j�  j  KbubKDj  )��}�(j�  KDj  ]�j�  j�  j  KbubKEj  )��}�(j�  KEj  ]�j�  j�  j  KbubKFj  )��}�(j�  KFj  ]�j�  j�  j  KbubKGj  )��}�(j�  KGj  ]�j�  j�  j  KbubKHj  )��}�(j�  KHj  ]�j�  j�  j  KbubKIj  )��}�(j�  KIj  ]�j�  j�  j  KbubKJj  )��}�(j�  KJj  ]�j�  j�  j  KbubKKj  )��}�(j�  KKj  ]�j�  j�  j  KbubKLj  )��}�(j�  KLj  ]�j�  j�  j  KbubKMj  )��}�(j�  KMj  ]�j�  j�  j  KbubKNj  )��}�(j�  KNj  ]�j�  j�  j  KbubKOj  )��}�(j�  KOj  ]�j�  j�  j  KbubKPj  )��}�(j�  KPj  ]�j�  j�  j  KbubKQj  )��}�(j�  KQj  ]�j�  j�  j  KbubKRj  )��}�(j�  KRj  ]�j�  j�  j  KbubKSj  )��}�(j�  KSj  ]�j�  j�  j  KbubKTj  )��}�(j�  KTj  ]�j�  j�  j  KbubKUj  )��}�(j�  KUj  ]�j�  j�  j  KbubKVj  )��}�(j�  KVj  ]�j�  j�  j  KbubKWj  )��}�(j�  KWj  ]�j�  j�  j  KbubKXj  )��}�(j�  KXj  ]�j�  j�  j  KbubKYj  )��}�(j�  KYj  ]�j�  j�  j  KbubKZj  )��}�(j�  KZj  ]�j�  j�  j  KbubK[j  )��}�(j�  K[j  ]�j�  j�  j  KbubK\j  )��}�(j�  K\j  ]�j�  j�  j  KbubK]j  )��}�(j�  K]j  ]�j�  j�  j  KbubK^j  )��}�(j�  K^j  ]�j�  j�  j  KbubK_j  )��}�(j�  K_j  ]�j�  j�  j  KbubK`j  )��}�(j�  K`j  ]�j�  j�  j  KbubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KbubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KbubKcj  )��}�(j�  Kcj  ]�j�  j�  j  KbubuKc}�(K j  )��}�(j�  K j  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubK	j  )��}�(j�  K	j  ]�j�  j�  j  KcubK
j  )��}�(j�  K
j  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubKj  )��}�(j�  Kj  ]�j�  j�  j  KcubK j  )��}�(j�  K j  ]�j�  j�  j  KcubK!j  )��}�(j�  K!j  ]�j�  j�  j  KcubK"j  )��}�(j�  K"j  ]�j�  j�  j  KcubK#j  )��}�(j�  K#j  ]�j�  j�  j  KcubK$j  )��}�(j�  K$j  ]�j�  j�  j  KcubK%j  )��}�(j�  K%j  ]�j�  j�  j  KcubK&j  )��}�(j�  K&j  ]�j�  j�  j  KcubK'j  )��}�(j�  K'j  ]�j�  j�  j  KcubK(j  )��}�(j�  K(j  ]�j�  j�  j  KcubK)j  )��}�(j�  K)j  ]�j�  j�  j  KcubK*j  )��}�(j�  K*j  ]�j�  j�  j  KcubK+j  )��}�(j�  K+j  ]�j�  j�  j  KcubK,j  )��}�(j�  K,j  ]�j�  j�  j  KcubK-j  )��}�(j�  K-j  ]�j�  j�  j  KcubK.j  )��}�(j�  K.j  ]�j�  j�  j  KcubK/j  )��}�(j�  K/j  ]�j�  j�  j  KcubK0j  )��}�(j�  K0j  ]�j�  j�  j  KcubK1j  )��}�(j�  K1j  ]�j�  j�  j  KcubK2j  )��}�(j�  K2j  ]�j�  j�  j  KcubK3j  )��}�(j�  K3j  ]�j�  j�  j  KcubK4j  )��}�(j�  K4j  ]�j�  j�  j  KcubK5j  )��}�(j�  K5j  ]�j�  j�  j  KcubK6j  )��}�(j�  K6j  ]�j�  j�  j  KcubK7j  )��}�(j�  K7j  ]�j�  j�  j  KcubK8j  )��}�(j�  K8j  ]�j�  j�  j  KcubK9j  )��}�(j�  K9j  ]�j�  j�  j  KcubK:j  )��}�(j�  K:j  ]�j�  j�  j  KcubK;j  )��}�(j�  K;j  ]�j�  j�  j  KcubK<j  )��}�(j�  K<j  ]�j�  j�  j  KcubK=j  )��}�(j�  K=j  ]�j�  j�  j  KcubK>j  )��}�(j�  K>j  ]�j�  j�  j  KcubK?j  )��}�(j�  K?j  ]�j�  j�  j  KcubK@j  )��}�(j�  K@j  ]�j�  j�  j  KcubKAj  )��}�(j�  KAj  ]�j�  j�  j  KcubKBj  )��}�(j�  KBj  ]�j�  j�  j  KcubKCj  )��}�(j�  KCj  ]�j�  j�  j  KcubKDj  )��}�(j�  KDj  ]�j�  j�  j  KcubKEj  )��}�(j�  KEj  ]�j�  j�  j  KcubKFj  )��}�(j�  KFj  ]�j�  j�  j  KcubKGj  )��}�(j�  KGj  ]�j�  j�  j  KcubKHj  )��}�(j�  KHj  ]�j�  j�  j  KcubKIj  )��}�(j�  KIj  ]�j�  j�  j  KcubKJj  )��}�(j�  KJj  ]�j�  j�  j  KcubKKj  )��}�(j�  KKj  ]�j�  j�  j  KcubKLj  )��}�(j�  KLj  ]�j�  j�  j  KcubKMj  )��}�(j�  KMj  ]�j�  j�  j  KcubKNj  )��}�(j�  KNj  ]�j�  j�  j  KcubKOj  )��}�(j�  KOj  ]�j�  j�  j  KcubKPj  )��}�(j�  KPj  ]�j�  j�  j  KcubKQj  )��}�(j�  KQj  ]�j�  j�  j  KcubKRj  )��}�(j�  KRj  ]�j�  j�  j  KcubKSj  )��}�(j�  KSj  ]�j�  j�  j  KcubKTj  )��}�(j�  KTj  ]�j�  j�  j  KcubKUj  )��}�(j�  KUj  ]�j�  j�  j  KcubKVj  )��}�(j�  KVj  ]�j�  j�  j  KcubKWj  )��}�(j�  KWj  ]�j�  j�  j  KcubKXj  )��}�(j�  KXj  ]�j�  j�  j  KcubKYj  )��}�(j�  KYj  ]�j�  j�  j  KcubKZj  )��}�(j�  KZj  ]�j�  j�  j  KcubK[j  )��}�(j�  K[j  ]�j�  j�  j  KcubK\j  )��}�(j�  K\j  ]�j�  j�  j  KcubK]j  )��}�(j�  K]j  ]�j�  j�  j  KcubK^j  )��}�(j�  K^j  ]�j�  j�  j  KcubK_j  )��}�(j�  K_j  ]�j�  j�  j  KcubK`j  )��}�(j�  K`j  ]�j�  j�  j  KcubKaj  )��}�(j�  Kaj  ]�j�  j�  j  KcubKbj  )��}�(j�  Kbj  ]�j�  j�  j  KcubKcj  )��}�(j�  Kcj  ]�j�  j�  j  Kcubuu�stairsUp�]�(K<K9e�SeenMap�]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKK K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKK K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K KKKK K KKKKKKKKK K K K K K K KKKK K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKK K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKK K K KKKK K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKK K K KKK K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K KKK K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKK K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K KKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K KKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKKKKK K K K K K K K K K K K K K K K K K KKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKKKKK K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKKKKK K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K KK K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKK K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKK K K K K K K K K K KKK K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKK K K K K K K K K K KKK K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K K K K K K K KKKKKKKKKKKKK K K K K KKKK K K K K K KKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K KKKKKKKKKKKK K KKKKKK K K K K KKKK K K K K K KKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKK K K K K K K K K K K K K K �       K K K K e]�(K KKKKKKKKKKKK K K K K K KKKKKKKKKKKK K KKKKKK K K K K KKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKK K K K K K KK K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K KKKK K K KKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK K K K K K KKKK K K KKKKKKKKKKKKK K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKK K KKKKK K K K K K KKKK K K KKKKKKKKKKKKK K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K KKKKKK K KKKKKKKKKKKKKK K K K KKKK K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K KKKKKK K KKKKKKKKKKKKKK K K K KKKK K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K KKKKKK K KKKKKKKKKKKKKK K K K KKKK K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K KKK K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K KKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K ee�djikstra_Player�j�  �master_Changed_Tiles�]�(]�(KCKe]�(KBKe]�(K>Ke]�(K?Ke]�(K?Ke]�(K>Ke]�(KQKDe]�(KQKFe]�(KQKDe]�(KQKFe]�(KQKDe]�(KQKFe]�(KQKDe]�(KQKFe]�(KQKDe]�(KQKFe]�(KQKDe]�(KQKFe]�(KQKDe]�(KRKFe]�(KQKGe]�(KQKHe]�(KPKIe]�(KPKJe]�(KOKKe]�(KOKLe]�(KNKMe]�(KRKDe]�(KQKCe]�(KRKFe]�(KQKGe]�(KQKHe]�(KPKIe]�(KPKJe]�(KPKKe]�(KOKLe]�(KOKMe]�(KRKDe]�(KQKCe]�(KRKFe]�(KQKGe]�(KQKHe]�(KQKIe]�(KPKJe]�(KPKKe]�(KPKLe]�(KOKMe]�(KRKDe]�(KQKCe]�(KRKFe]�(KRKGe]�(KQKHe]�(KQKIe]�(KQKJe]�(KQKKe]�(KPKLe]�(KPKMe]�(KRKDe]�(KRKCe]�(KQKBe]�(KRKFe]�(KRKGe]�(KRKHe]�(KQKIe]�(KQKJe]�(KQKKe]�(KQKLe]�(KQKMe]�(KRKDe]�(KRKCe]�(KRKBe]�(KRKAe]�(KRK@e]�(KQK?e]�(KQK>e]�(KQK=e]�(KRKFe]�(KRKGe]�(KRKHe]�(KRKIe]�(KRKJe]�(KRKKe]�(KQKLe]�(KQKMe]�(KRKDe]�(KRKCe]�(KRKBe]�(KRKAe]�(KRK@e]�(KRK?e]�(KRKFe]�(KRKGe]�(KRKHe]�(KRKIe]�(KRKJe]�(KRKKe]�(KRKLe]�(KRKMe]�(KRKDe]�(KRKCe]�(KRKBe]�(KRKAe]�(KRK@e]�(KSK?e]�(KRKFe]�(KRKGe]�(KRKHe]�(KRKIe]�(KRKJe]�(KRKKe]�(KSKLe]�(KSKMe]�(KRKDe]�(KRKCe]�(KSKBe]�(KRKFe]�(KRKGe]�(KRKHe]�(KSKIe]�(KSKJe]�(KSKKe]�(KSKLe]�(KSKMe]�(KRKDe]�(KSKCe]�(KRKFe]�(KRKGe]�(KSKHe]�(KSKIe]�(KSKJe]�(KSKKe]�(KTKLe]�(KTKMe]�(KRKDe]�(KSKCe]�(KRKFe]�(KSKGe]�(KSKHe]�(KSKIe]�(KTKJe]�(KTKKe]�(KTKLe]�(KUKMe]�(KRKDe]�(KSKCe]�(KRKFe]�(KSKGe]�(KSKHe]�(KTKIe]�(KTKJe]�(KTKKe]�(KUKLe]�(KSKDe]�(KRKFe]�(KSKGe]�(KSKHe]�(KTKIe]�(KTKJe]�(KUKKe]�(KSKDe]�(KSKFe]�(KSKDe]�(KSKFe]�(KSKDe]�(KSKFe]�(KSKDe]�(KSKFe]�(KSKDe]�(KSKFe]�(KSKDe]�(KSKFe]�(KQKDe]�(KSKDe]�(KQKDe]�(KSKDe]�(KQKDe]�(KSKDe]�(KQKDe]�(KSKDe]�(KQKDe]�(KSKDe]�(KQKDe]�(KSKDe]�(KQKDe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKEe]�(KSKEe]�(KQKFe]�(KSKEe]�(KQKFe]�(KSKFe]�(KQKFe]�(KSKFe]�(KQKFe]�(KSKFe]�(KQKFe]�(KSKFe]�(KQKFe]�(KSKFe]�(KQKFe]�(KSKFeej�  h�SeesMap�]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K ee�CollisionMap�]�(]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K KKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K KKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKK KKKKKKKKKKKKKKKKKKKK KKKKKK K K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKK KKKKKKKKKKKKKKKKKKKK KKKKKK K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKK KKKKK K K K K K KKKKKKKKKK KKKKKK KKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K KKKKKK KKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKKKKKKK K K K KKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKKKKKKK K K K KKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K KKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKK K K KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K KKKKKKKKKKKK KKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKK KKKKKKKKKKKK KKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKKKKKKKK K K KKKKK K K KKKKKKKK KKKKKKKKKKKK KKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKKKKKKKK K K KKKKK K K KKKKKKKK KKKKKKKKK K K K K K K K K KKKKKKKKK K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK K K K K K K K K KKKKK K K KKKKKKKK KKKKKKKKK K K K K K K K K KKKKKKKKK KKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K KKKKK K K KKKKKKKK K K K K K K K K K K K K K K K K K KKKKKKKKK KKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKK KKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K KKKKK K KKKKKKKKK KKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKK KKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K KKKKK K KKKKKKKKK KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKK KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K KKKKK K KKKKKKKKK KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K KKKKK K K K K K K K K K K KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K K KKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKK K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKe]�(KKK K K KKK K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKe]�(KKK K K KKK K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K KKKKKKKKK KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKK K K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K K K K K K K K K KKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K KKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKK KKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKK KKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K KKKKKKKK KKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKK KKKKKKKK KKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K KKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKK KKKKKKKK KKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKK KKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKK KKKKKKKK K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKK K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKK K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK K K K KKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK KKKKKKKKKKKKKKKKKKKKKKKKKK K K KKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK KKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K K K K K KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K KKKKK KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKK K KKKK K K KKKKK KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKK K KKKK K K KKKKK KKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKK K KKKK K K KKKKK KKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K KKKKK KKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K KKK K K KKKKKKKKK KKKKKKKK K K K K K K K KKKKK KKKKKKKKK K K K K K K K K K K K K K K K K K K KKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K KKK K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKK KKKKKKKKK K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKee�itemList�]�(jf  j
  j  h�h�h7�Staff���j  h7�Buckler���hzhshOh�hjh�h�hhbhZhX�Iron_Breastplate���hnh�j  eh^j�  �djikstra_Player_Adj�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNKOKPKQNNNNNNNNNNNNNNNNNK[K\K]K^K_K`NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKpKoKnKmKlKkKjNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKMKNKOKPNNNNNNNNNNNNNNNNNKZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKoKnKmKlKkKjKiNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKJKKKLKMKNKONNNNNNNNNNNNNNNNNKYKZK[K\K]K^NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKnKmKlKkKjKiKhKgKfKeKdKcKbKaK`K_NNNNNNNNNNNNNNNNNNNKOKNKMKLKKKJKIKJKKKLKMKNNNNNNNNNNNNNNNNNNKXKYKZK[K\K]K^K_K`NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKoKnKmKlKkKjKiNNNNNNNNK^NNNNNNNNNNNNNNNNNNNKPNNNNNKHKIKJKKKLKMNNNNNNNNNNNNNNNNNKWKXKYKZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKpKoKnKmKlKkKjNNNNNNNNK]NNNNNNNNNNNNNNNNNNNKQNNNNNKGKHKIKJKKKLKMKNKOKPKQKRKSKTKUKVNNNNNNNKVKWKXKYKZK[K\K]K^NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKqKpKoKnKmKlKkNNNNNNNNK\NNNNKWKVKUKTKUKVNNNNNNNNNKRNNNNNKFNNNNNNNNNNNNNNKWKXKYKZKYKXKWKVKUKVKWKXKYKZK[K\K]NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKrKqKpKoKnKmKlNNNNNNNNK[KZKYKXKWKVKUKTKSKTKUKVKWKXKYKXKWKVKUKTKSNNNNNKENNNNNNNNNNNNNNNNNNNNNNKTKUKVKWKXKYKZK[K\NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKsKrKqKpKoKnKmNNNNNNNNNNNNNKUKTKSKRNNNNNNNNNNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNNNKSNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKtKsKrKqKpKoKnNNNNNNNNNNNNNKTKSKRKQNNNNNNNNNNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNNNKRNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKuKtKsKrKqKpKoNNNNNNNNNNNNNKSKRKQKPKQKRNNNNNNNNNNNNNNNKBNNNNNNNNNNNNNNNNNNNNNNKQNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKtNNNNNNNNNNNNNNNNNKRKQKPKOKPKQNNNNNNNNNNNNNNNKANNNNNNNNNNNNNNNNNNNNNNKPNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKuNNNNNNNNNNNNNNNNNKQKPKOKNKOKPNNNNNNNNNNNNNNNK@NNNNNNNNNNNNNNNNNNNNNNKONNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKvNNNNNNNNNNNNNNNNNKPKOKNKMKNKONNNNNNNNNNNNNNNK?NNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKwNNNNNNNNNNNNNNNNNNNNKLNNNNNNNNNNNNNNNNNK>K=K<K;K:K9K8NNNNNNNNNNNNNNNNKMNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKxNNNNNNNNNNNNNNNNNNNNKKNNNNNNNNNNNNNNNNNNNNNNNK7NNNNNNNNNNNNNNNNKLNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKyNNNNNNNNNNNNNNNNNNNNKJNNNNNNNNNNNNNNNNNNNNNNNK6NNNNNNNNNNNNNNNNKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKxNNNNNNNNNNNNNNNNNNNNKIKHNNNNNNNNNNNNNNNNNNNNNNK5NNNNNNNNNNNNNNNNKJKIKHNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKwNNNNNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKsKtKuKvNNNNNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKrNNNNNNNNNNNNNNNNNNKKKJKIKHKGKFKEKDKCKBNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNKENNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKqNNNNNNNNNNNNNNNNNNKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKpNNNNNNNNNNNNNNNNNNKKKJKIKHKGKFKEKDKCKBNNNNNNNK8NNNNNNNNNNNK0NNNNNNNNNNNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqKpKoKnKmKlKkNNNNNNNNNNNNNNKLKKKJNNNNKEKDKCNNNNNNNK7NNNNNNNNNNNK/NNNNNNNNNNNNNNNNK@KAKBKCKBKCKDKEKFKGNNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpKoKnKmKlKkKjNNNNNNNNNNNNNNKMKLKKNNNNKFKEKDNNNNNNNK6NNNNNNNNK-K,K-K.K/K0K1K2K3NNNNNNNNK<K=K>K?K@KAKBKAKBKCKDKEKFNNNNNNNNNNNNNNNNNNNe]�(NNKqKpKoKnKmKlKkKjKiNNNNNNNNKTKSKRKQKPKOKNKMKLNNNNKGKFKENNNNNNNK5NNNNNNNNK,K+K,K-K.K/K0K1K2NNNNNNNNK;NNK@KAKBKAK@KAKBKCKDKENNNNNNNNNNNNNNNNNNNe]�(NNKpKoKnKmKlKkKjKiKhNNNNNNNNKUNNNNNKOKNKMNNNNKHKGKFNNNNNNNK4K3K2K1K0K/K.K-K,K+K*K+K,K-K.K/K0K1NNNNNNNNK:NNKAKBKAK@K?K@KAKBKCKDNNNNNNNNNNNNNNNNNNNe]�(NNKoKnKmKlKkKjKiKhKgNNNNNNNNKVNNNNNKPKOKNKMKLKKKJKIKHKGNNNNNNNNNNNNNNNNK*K)K*K+K,K-K.K/K0NNNNNNNNK9NNNNK@K?K>K?K@KAKBKCNNNNNNNNNNNNNNNNNNNe]�(NNKpKoKnNNNNKgKfNNNNNNNNKWNNNNNKQKPKOKNKMKLKKKJKIKHNNNNNNNNNNNNNNNNK)K(K)K*K+K,K-K.K/NNNNNNNNK8NNNNK?K>K=K>K?K@KAKBNNNNNNNNNNNNNNNNNNNe]�(NNKqKpKoNNNNKfKeNNNNNNNNKXNNNNNNKQNNNNNNNNNNNNNNNNNNNNNNNNK(K'K(K)K*K+K,K-K.NNNNNNNNK7NNNNNNK<NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpNNNNKeKdNNNNNNNNKYNNNNNNKRNNNNNNNNNNNNNNNNNNNNNNNNK'K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6NNNNNNK;NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqNNNNKdKcKbKaK`K_K^K]K\K[KZNNNNNNKSNNNNNNNNNNNNNNNNNNNNNNNNNK%NNNNNNNNNNNNNNNNNNNNNNK:K9K8K7K6NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKeNNNNNNNNNNNNNNNNKTNNNNNNNNNNNNNNNNNNNNNNNNNK$NNNNNNNNNNNNNNNNNNNNNNNNNNK5NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKfNNNNNNNNNNNNNNNNKUNNNNNNNNNNNNNNNNNNNNNNNNNK#K"K!K KNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKgNNNNNNNNNNNNNNNNKVNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNe]�(NNNNKmKlKkKjKiKhNNNNNNNNNNNNNNNNKWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNe]�(NNNNKnNNNNNNNNNNNNNNNNNNNNNKXNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNe]�(NNNNKoNNNNNNNNNNNNNNNNNNNNNKYNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNK0K1K0K/K0NNNNNNNNNNNNNNNNNNe]�(NNNNKpNNNNNNNNNNNNNNNNNNNNNKZNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNK/K0K/K.K/NNNNNNNNNNNNNNNNNNe]�(NNNNKqNNNNNNNNNNNNNNNNNNNNNK[NNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNK.K/K.K-K.NNNNNNNNNNNNNNNNNNe]�(NNNNKrNNNNNNNNNNNNNNNNNNNNK]K\K]K^K_K`KaKbKcNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNK*K+K,K-K.K-K,K-NNNNNNNNNNNNNNNNNNe]�(NNNNKsNNNNNNNNNNNNNNKdKcKbKaK`K_K^K]K^K_K`KaKbKcKdNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNK)K*K+K,K-K,K+K,NNNNNNNNNNNNNNNNNNe]�(NNKvKuKtKuKvKwKxKyKzNNNNNNNNKeNNNNNK_K^K_K`KaKbKcKdKeNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNK"K#K$K%K&K'K(K)K*K+K,K+K*K+NNNNNNNNNNNNNNNNNNe]�(NNKwKvKuKvKwKxKyKzK{NNNNNNNNKfNNNNNK`K_K`K_K`KaKbKcKdNNNNNNNNNNNNNNNNKKKKKKKKKKKKKKKKKK K!NNNNNK)K*K+K,K+K*K)K*NNNNNNNNNNNNNNNNNNe]�(NNKvKuKtKuKvKwKxKyKzNNNNNNNNKgNNNNNKaK`K_K^K_K`KaKbKcNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNK*K+K,K+K*K)K(K)NNNNNNNNNNNNNNNNNNe]�(NNKuKtKsNNKvKwKxKyNNNNNNNNKhNNNNNK`K_K^K]K^K_K`KaKbNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNK'NNNNNNNNNNNNNNNNNNNe]�(NNKtKsKrNNKuKvKwKxNNNNNNNNKiNNNNNK_K^K]K\K]K^K_K`KaNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNK&NNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqKrKsKtKuKvKwNNNNNNNNKjNNNNNK^K]K\K[K\K]K^K_K`NNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNK%NNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpKqKrKsKtKuKvNNNNNNNNKkNNNNNK]K\K[KZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNKKKKKKK K!K"K#K$NNNNNNNNNNNNNNNNNNNe]�(NNKqKpKoKpKqKrKsKtKuKtKsKrKqKpKoKnKmKlNNNNNK\K[KZKYKZK[K\K]K^NNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKnNNNNNNNNNNNNNNNNNNNNNNNKXNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKmKlKkKjKiNNNNNNNNNNNNNNNNNNNKWNNNNNNNNNNNNNNNNNNNNNNNNNKK
K	KKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKhNNNNNNNNNNNNNNNNNNNKVNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKgNNNNNNNNNNNNNNNNNNNKUKTKSKRKQNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKlKkKjKiKhKgKfKeKdKcNNNNNNNNNNNNNNNNNNNNKPNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKkKjKiKhKgKfKeKdKcKbNNNNNNNNNNNNNNNNNNNNKONNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKjKiKhKgKfKeKdKcKbKaK`K_K^K]K\K[KZKYNNNNNNNNNKOKNKMKNKONNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKkKjKiKhKgKfKeKdKcKbNNNNNNNKXNNNNNNNNNKNKMKLKMKNNNNNNNNNNNNNNNNNNNKKKKKK KNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKlKkKjKiKhKgNNNKcNNNNNNNKWNNNNNNNKOKNKMKLKKKLKMNNNNNNNNNNNNNNNNNNKKKKK KK KKKKKKKKNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKmKlKkKjKiKhNNNKdNNNNNNNKVNNNNNNNKNKMKLKKKJKKKLNNNNNNNNNNNNNNNNNNKKKKKK KNNNNNNNK	NNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKnKmKlKkKjKiNNNKeNNNNNNNKUKTKSKRKQKPKOKNKMKLKKKJKIKJKKNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNK
KKKKKKKKKKKNNNNNNNNNN�      NNNNNNNNNNNNe]�(NNKoKnKmKlKkKjKiKhKgKfNNNNNNNNNNNNNNNKLKKKJKIKHKIKJNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKlNNNNNNNNNNNNNNNNNNNNKKKJKIKHKGKHKINNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKmNNNNNNNNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNK	KKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKnNNNNNNNNNNNNNNNNNNNNNNNNKENNNNNNNNNNNNNNNNNNNNK
K	KKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKmNNNNNNNNNNNNNNNNNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNKK
K	KKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKlNNNNNNNNNNNNNNNNNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNKKK
K	KKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKhKiKjKkNNNNNNNNNNNNNNNNNNNNNNNNKBNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKgNNNNNNNNNNNNNNNNNNNNNNNNNNNKANNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKfNNNNNNNNNNNNNNNNNNNNNNNNNK>K?K@NNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKeNNNNNNNNNNNNNNNNNNNNNNNNNK=NNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKdNNNNNNNNNNNNNNNNNNNNNNNNNK<NNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKcNNNNNNNNNNNNNNNNNNNNNK?K>K=K<K;K:K9K8NNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKcKbKaK`K_K^K]NNNNNNNNNNNNNNNNK>K=K<K;K:K9K8K7K6K5K4K3K2NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKbKaK`K_K^K]K\NNNNNNNNNNNNNNNNK?K>K=K<K;K:K9K8NNNNK1NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKaK`K_K^K]K\K[NNNNNNNNNNNNNNNNK@K?NNNK;K:K9NNNNK0NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK`K_K^K]K\K[KZNNNNNNNNNNNNNNNNKAK@NNNK<K;K:NNNNK/NNNNNNNNKKKKKKK K!NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK_K^K]K\K[KZKYNNNNNNNNNNNNNNNNKBKANNNK=K<K;NNNNK.NNNNNNNNKKKKKK K!K"NNNNNNNNNNNNNNNNNK:K;K<K=K>K?K@KAKBKCNNNNNNNNNNNNNNNNNNNe]�(NNK^K]K\K[KZKYKXNNNNNNNNKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NNNNK-NNNNNNNNKKKKK K!K"K#NNNNNNNNNNNNNNNNNK9K:K;K<K=K>K?K@KAKBNNNNNNNNNNNNNNNNNNNe]�(NNK_K^NNKYKXKWNNNNNNNNKLNNNNNNNKDKCKBKAK@K?K>K=NNNNK,NNNNNNNNKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/NNNNNNK8K9K:K;K<K=K>K?K@KANNNNNNNNNNNNNNNNNNNe]�(NNK^K]NNKXKWKVKUKTKSKRKQKPKOKNKMNNNNNNNNNNNNNNNNNNNK+NNNNNNNNK KK K!K"K#K$K%NNNNNNNNNNK0K1K2K3K4K5K6K7K8K9K:K;K<K=K>K?K@NNNNNNNNNNNNNNNNNNNe]�(NNK]K\K[KZKYKXKWNNNNNNNNNNNNNNNNNNNNNNNNNNNNK*K)K(K'K&K%K$K#K"K!K K!K"K#K$K%K&NNNNNNNNNNNNNNNNNK8K9K:K;K<K=K>K?K@KANNNNNNNNNNNNNNNNNNNe]�(NNK^K]K\K[KZKYKXNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK#K$K%K&K'NNNNNNNNNNNNNNNNNK9K:K;K<K=K>K?K@KAKBNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK$K%K&K'K(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK%K&K'K(K)NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej�  j�  �
stairsDown�]�(KSKOe�djikstra_Stairs_Up�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKOKPKQKRNNNNNNNNNNNNNNNNNK\K]K^K_K`KaNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKqKpKoKnKmKlKkNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNKOKPKQNNNNNNNNNNNNNNNNNK[K\K]K^K_K`NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKpKoKnKmKlKkKjNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKLKMKNKOKPNNNNNNNNNNNNNNNNNKZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKoKnKmKlKkKjKiKhKgKfKeKdKcKbKaK`NNNNNNNNNNNNNNNNNNNKPKOKNKMKLKKKJKKKLKMKNKONNNNNNNNNNNNNNNNNKYKZK[K\K]K^K_K`KaNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKpKoKnKmKlKkKjNNNNNNNNK_NNNNNNNNNNNNNNNNNNNKQNNNNNKIKJKKKLKMKNNNNNNNNNNNNNNNNNNKXKYKZK[K\K]K^K_K`NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKqKpKoKnKmKlKkNNNNNNNNK^NNNNNNNNNNNNNNNNNNNKRNNNNNKHKIKJKKKLKMKNKOKPKQKRKSKTKUKVKWNNNNNNNKWKXKYKZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKrKqKpKoKnKmKlNNNNNNNNK]NNNNKXKWKVKUKVKWNNNNNNNNNKSNNNNNKGNNNNNNNNNNNNNNKXKYKZK[KZKYKXKWKVKWKXKYKZK[K\K]K^NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKsKrKqKpKoKnKmNNNNNNNNK\K[KZKYKXKWKVKUKTKUKVKWKXKYKZKYKXKWKVKUKTNNNNNKFNNNNNNNNNNNNNNNNNNNNNNKUKVKWKXKYKZK[K\K]NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKtKsKrKqKpKoKnNNNNNNNNNNNNNKVKUKTKSNNNNNNNNNNNNNNNNNKENNNNNNNNNNNNNNNNNNNNNNKTNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKuKtKsKrKqKpKoNNNNNNNNNNNNNKUKTKSKRNNNNNNNNNNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNNNKSNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKvKuKtKsKrKqKpNNNNNNNNNNNNNKTKSKRKQKRKSNNNNNNNNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNNNKRNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKuNNNNNNNNNNNNNNNNNKSKRKQKPKQKRNNNNNNNNNNNNNNNKBNNNNNNNNNNNNNNNNNNNNNNKQNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKvNNNNNNNNNNNNNNNNNKRKQKPKOKPKQNNNNNNNNNNNNNNNKANNNNNNNNNNNNNNNNNNNNNNKPNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKwNNNNNNNNNNNNNNNNNKQKPKOKNKOKPNNNNNNNNNNNNNNNK@NNNNNNNNNNNNNNNNNNNNNNKONNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKxNNNNNNNNNNNNNNNNNNNNKMNNNNNNNNNNNNNNNNNK?K>K=K<K;K:K9NNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKyNNNNNNNNNNNNNNNNNNNNKLNNNNNNNNNNNNNNNNNNNNNNNK8NNNNNNNNNNNNNNNNKMNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKzNNNNNNNNNNNNNNNNNNNNKKNNNNNNNNNNNNNNNNNNNNNNNK7NNNNNNNNNNNNNNNNKLNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKyNNNNNNNNNNNNNNNNNNNNKJKINNNNNNNNNNNNNNNNNNNNNNK6NNNNNNNNNNNNNNNNKKKJKINNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKxNNNNNNNNNNNNNNNNNNNNNKHNNNNNNNNNNNNNNNNNNNNNNK5NNNNNNNNNNNNNNNNNNKHNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKtKuKvKwNNNNNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKsNNNNNNNNNNNNNNNNNNKLKKKJKIKHKGKFKEKDKCNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKrNNNNNNNNNNNNNNNNNNKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNKENNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKqNNNNNNNNNNNNNNNNNNKLKKKJKIKHKGKFKEKDKCNNNNNNNK9NNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKtKsKrKqKpKoKnKmKlNNNNNNNNNNNNNNKMKLKKNNNNKFKEKDNNNNNNNK8NNNNNNNNNNNK0NNNNNNNNNNNNNNNNKAKBKCKDKCKDKEKFKGKHNNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqKpKoKnKmKlKkNNNNNNNNNNNNNNKNKMKLNNNNKGKFKENNNNNNNK7NNNNNNNNK.K-K.K/K0K1K2K3K4NNNNNNNNK=K>K?K@KAKBKCKBKCKDKEKFKGNNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpKoKnKmKlKkKjNNNNNNNNKUKTKSKRKQKPKOKNKMNNNNKHKGKFNNNNNNNK6NNNNNNNNK-K,K-K.K/K0K1K2K3NNNNNNNNK<NNKAKBKCKBKAKBKCKDKEKFNNNNNNNNNNNNNNNNNNNe]�(NNKqKpKoKnKmKlKkKjKiNNNNNNNNKVNNNNNKPKOKNNNNNKIKHKGNNNNNNNK5K4K3K2K1K0K/K.K-K,K+K,K-K.K/K0K1K2NNNNNNNNK;NNKBKCKBKAK@KAKBKCKDKENNNNNNNNNNNNNNNNNNNe]�(NNKpKoKnKmKlKkKjKiKhNNNNNNNNKWNNNNNKQKPKOKNKMKLKKKJKIKHNNNNNNNNNNNNNNNNK+K*K+K,K-K.K/K0K1NNNNNNNNK:NNNNKAK@K?K@KAKBKCKDNNNNNNNNNNNNNNNNNNNe]�(NNKqKpKoNNNNKhKgNNNNNNNNKXNNNNNKRKQKPKOKNKMKLKKKJKINNNNNNNNNNNNNNNNK*K)K*K+K,K-K.K/K0NNNNNNNNK9NNNNK@K?K>K?K@KAKBKCNNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpNNNNKgKfNNNNNNNNKYNNNNNNKRNNNNNNNNNNNNNNNNNNNNNNNNK)K(K)K*K+K,K-K.K/NNNNNNNNK8NNNNNNK=NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqNNNNKfKeNNNNNNNNKZNNNNNNKSNNNNNNNNNNNNNNNNNNNNNNNNK(K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7NNNNNNK<NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKtKsKrNNNNKeKdKcKbKaK`K_K^K]K\K[NNNNNNKTNNNNNNNNNNNNNNNNNNNNNNNNNK&NNNNNNNNNNNNNNNNNNNNNNK;K:K9K8K7NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKfNNNNNNNNNNNNNNNNKUNNNNNNNNNNNNNNNNNNNNNNNNNK%NNNNNNNNNNNNNNNNNNNNNNNNNNK6NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKgNNNNNNNNNNNNNNNNKVNNNNNNNNNNNNNNNNNNNNNNNNNK$K#K"K!K NNNNNNNNNNNNNNNNNNNNNNK5NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKhNNNNNNNNNNNNNNNNKWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNNNe]�(NNNNKnKmKlKkKjKiNNNNNNNNNNNNNNNNKXNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNe]�(NNNNKoNNNNNNNNNNNNNNNNNNNNNKYNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNe]�(NNNNKpNNNNNNNNNNNNNNNNNNNNNKZNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNK1K2K1K0K1NNNNNNNNNNNNNNNNNNe]�(NNNNKqNNNNNNNNNNNNNNNNNNNNNK[NNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNK0K1K0K/K0NNNNNNNNNNNNNNNNNNe]�(NNNNKrNNNNNNNNNNNNNNNNNNNNNK\NNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNK/K0K/K.K/NNNNNNNNNNNNNNNNNNe]�(NNNNKsNNNNNNNNNNNNNNNNNNNNK^K]K^K_K`KaKbKcKdNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNK+K,K-K.K/K.K-K.NNNNNNNNNNNNNNNNNNe]�(NNNNKtNNNNNNNNNNNNNNKeKdKcKbKaK`K_K^K_K`KaKbKcKdKeNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNK*K+K,K-K.K-K,K-NNNNNNNNNNNNNNNNNNe]�(NNKwKvKuKvKwKxKyKzK{NNNNNNNNKfNNNNNK`K_K`KaKbKcKdKeKfNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNK#K$K%K&K'K(K)K*K+K,K-K,K+K,NNNNNNNNNNNNNNNNNNe]�(NNKxKwKvKwKxKyKzK{K|NNNNNNNNKgNNNNNKaK`KaK`KaKbKcKdKeNNNNNNNNNNNNNNNNKKKKKKKKKKKKKKKKK K!K"NNNNNK*K+K,K-K,K+K*K+NNNNNNNNNNNNNNNNNNe]�(NNKwKvKuKvKwKxKyKzK{NNNNNNNNKhNNNNNKbKaK`K_K`KaKbKcKdNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNK+K,K-K,K+K*K)K*NNNNNNNNNNNNNNNNNNe]�(NNKvKuKtNNKwKxKyKzNNNNNNNNKiNNNNNKaK`K_K^K_K`KaKbKcNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNK(NNNNNNNNNNNNNNNNNNNe]�(NNKuKtKsNNKvKwKxKyNNNNNNNNKjNNNNNK`K_K^K]K^K_K`KaKbNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNK'NNNNNNNNNNNNNNNNNNNe]�(NNKtKsKrKsKtKuKvKwKxNNNNNNNNKkNNNNNK_K^K]K\K]K^K_K`KaNNNNNNNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNK&NNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqKrKsKtKuKvKwNNNNNNNNKlNNNNNK^K]K\K[K\K]K^K_K`NNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNKKKKKK K!K"K#K$K%NNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpKqKrKsKtKuKvKuKtKsKrKqKpKoKnKmNNNNNK]K\K[KZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKoNNNNNNNNNNNNNNNNNNNNNNNKYNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKnKmKlKkKjNNNNNNNNNNNNNNNNNNNKXNNNNNNNNNNNNNNNNNNNNNNNNNKKK
K	KNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKiNNNNNNNNNNNNNNNNNNNKWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKhNNNNNNNNNNNNNNNNNNNKVKUKTKSKRNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKmKlKkKjKiKhKgKfKeKdNNNNNNNNNNNNNNNNNNNNKQNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKlKkKjKiKhKgKfKeKdKcNNNNNNNNNNNNNNNNNNNNKPNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKkKjKiKhKgKfKeKdKcKbKaK`K_K^K]K\K[KZNNNNNNNNNKPKOKNKOKPNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKlKkKjKiKhKgKfKeKdKcNNNNNNNKYNNNNNNNNNKOKNKMKNKONNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKmKlKkKjKiKhNNNKdNNNNNNNKXNNNNNNNKPKOKNKMKLKMKNNNNNNNNNNNNNNNNNNNKKKKKK KKKKKKKKK	NNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKnKmKlKkKjKiNNNKeNNNNNNNKWNNNNNNNKOKNKMKLKKKLKMNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNK
NNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKoKnKmKlKkKjNNNKfNNNNNNNKVKUKTKSKRKQKPKOKNKMKLKKKJKKKLNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNKKKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNKpKoKnKmKlKkKjKiKhKgNNNNNNNNNNNNNNNKMKLKKKJKIKJKKNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKmNNNNNNNNNNNNNNNNNNNNKLKKKJKIKHKIKJNNNNNNNNNNNNNNNNNNK	KKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKnNNNNNNNNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNK
K	KKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKoNNNNNNNNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNKK
K	KKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKnNNNNNNNNNNNNNNNNNNNNNNNNKENNNNNNNNNNNNNNNNNNNNKKK
K	KKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKmNNNNNNNNNNNNNNNNNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNKKKK
K	KK	NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKiKjKkKlNNNNNNNNNNNNNNNNNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKhNNNNNNNNNNNNNNNNNNNNNNNNNNNKBNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKgNNNNNNNNNNNNNNNNNNNNNNNNNK?K@KANNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKfNNNNNNNNNNNNNNNNNNNNNNNNNK>NNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKeNNNNNNNNNNNNNNNNNNNNNNNNNK=NNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKdNNNNNNNNNNNNNNNNNNNNNK@K?K>K=K<K;K:K9NNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKdKcKbKaK`K_K^NNNNNNNNNNNNNNNNK?K>K=K<K;K:K9K8K7K6K5K4K3NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKcKbKaK`K_K^K]NNNNNNNNNNNNNNNNK@K?K>K=K<K;K:K9NNNNK2NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKbKaK`K_K^K]K\NNNNNNNNNNNNNNNNKAK@NNNK<K;K:NNNNK1NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKaK`K_K^K]K\K[NNNNNNNNNNNNNNNNKBKANNNK=K<K;NNNNK0NNNNNNNNKKKKKK K!K"NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK`K_K^K]K\K[KZNNNNNNNNNNNNNNNNKCKBNNNK>K=K<NNNNK/NNNNNNNNKKKKK K!K"K#NNNNNNNNNNNNNNNNNK;K<K=K>K?K@KAKBKCKDNNNNNNNNNNNNNNNNNNNe]�(NNK_K^K]K\K[KZKYNNNNNNNNKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=NNNNK.NNNNNNNNKKKK K!K"K#K$NNNNNNNNNNNNNNNNNK:K;K<K=K>K?K@KAKBKCNNNNNNNNNNNNNNNNNNNe]�(NNK`K_NNKZKYKXNNNNNNNNKMNNNNNNNKEKDKCKBKAK@K?K>NNNNK-NNNNNNNNK KK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0NNNNNNK9K:K;K<K=K>K?K@KAKBNNNNNNNNNNNNNNNNNNNe]�(NNK_K^NNKYKXKWKVKUKTKSKRKQKPKOKNNNNNNNNNNNNNNNNNNNNK,NNNNNNNNK!K K!K"K#K$K%K&NNNNNNNNNNK1K2K3K4K5K6K7K8K9K:K;K<K=K>K?K@KANNNNNNNNNNNNNNNNNNNe]�(NNK^K]K\K[KZKYKXNNNNNNNNNNNNNNNNNNNNNNNNNNNNK+K*K)K(K'K&K%K$K#K"K!K"K#K$K%K&K'NNNNNNNNNNNNNNNNNK9K:K;K<K=K>K?K@KAKBNNNNNNNNNNNNNNNNNNNe]�(NNK_K^K]K\K[KZKYNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK$K%K&K'K(NNNNNNNNNNNNNNNNNK:K;K<K=K>K?K@KAKBKCNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK%K&K'K(K)NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK&K'K(K)K*NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�maze�]�(]�(�#�j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  �.�j�}  j�}  �x�j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  �=�j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  hCj�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  ji  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  �~�j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  ji  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  hCj�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  ji  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  hCj�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  �S�j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  hCj�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  �E�j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  hCj�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  �      j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  e]�(j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  j�}  ee�	enemyList�]�(�Enemies.Goblins��Goblin_Stonewall���j ~  �Goblin_Lancer���j ~  �Goblin_Berserker���j ~  �Goblin_Archer���j ~  �Goblin_Knight���j ~  �Goblin_Grunt���j ~  �Goblin_Thief���e�djikstra_Stairs_Down�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK�K�K�K�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK�K�K�K�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNK�K�K�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNK�NNNNNNNNNNNNNNNNNNNK�NNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNK�NNNNNNNNNNNNNNNNNNNK�NNNNNK�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�NNNNNNNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNK�NNNNK�K�K�K�K�K�NNNNNNNNNK�NNNNNK�NNNNNNNNNNNNNNK�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNK�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�NNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNK�K�K�K�NNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNK�K�K�K�NNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNK�KK~K}K|K{KzNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNKyNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNKxNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNK�K�NNNNNNNNNNNNNNNNNNNNNNKwNNNNNNNNNNNNNNNNK�K�K�NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNKvNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�K�K�K�NNNNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNKuNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNK}K|K}K~KK�K�K�K�K�NNNNNNNNNNNNNNNNNNNKtNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNK|K{K|K}K~KK�K�K�K�K�K�K�KK~K}K|K{NNNNNNNNNNNKsNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNK{KzK{K|K}K~KK�K�K�NNNNNNNKzNNNNNNNNNNNKrNNNNNNNNNNNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNKzKyKzNNNNKK�K�NNNNNNNKyNNNNNNNNNNNKqNNNNNNNNNNNNNNNNK�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNKyKxKyNNNNK~KK�NNNNNNNKxNNNNNNNNKoKnKoKpKqKrKsKtKuNNNNNNNNK~KK�K�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK~K}K|K{KzKyKxKwKxNNNNK}K~KNNNNNNNKwNNNNNNNNKnKmKnKoKpKqKrKsKtNNNNNNNNK}NNK�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNKNNNNNKwKvKwNNNNK|K}K~NNNNNNNKvKuKtKsKrKqKpKoKnKmKlKmKnKoKpKqKrKsNNNNNNNNK|NNK�K�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK�NNNNNKvKuKvKwKxKyKzK{K|K}NNNNNNNNNNNNNNNNKlKkKlKmKnKoKpKqKrNNNNNNNNK{NNNNK�K�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK�K�NNNNNNNNK�NNNNNKuKtKuKvKwKxKyKzK{K|NNNNNNNNNNNNNNNNKkKjKkKlKmKnKoKpKqNNNNNNNNKzNNNNK�K�KK�K�K�K�K�NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK�K�NNNNNNNNK�NNNNNNKsNNNNNNNNNNNNNNNNNNNNNNNNKjKiKjKkKlKmKnKoKpNNNNNNNNKyNNNNNNK~NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK�K�NNNNNNNNK�NNNNNNKrNNNNNNNNNNNNNNNNNNNNNNNNKiKhKiKjKkKlKmKnKoKpKqKrKsKtKuKvKwKxNNNNNNK}NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK�K�K�K�K�K�K�K�K�K�K�NNNNNNKqNNNNNNNNNNNNNNNNNNNNNNNNNKgNNNNNNNNNNNNNNNNNNNNNNK|K{KzKyKxNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNKpNNNNNNNNNNNNNNNNNNNNNNNNNKfNNNNNNNNNNNNNNNNNNNNNNNNNNKwNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNKoNNNNNNNNNNNNNNNNNNNNNNNNNKeKdKcKbKaNNNNNNNNNNNNNNNNNNNNNNKvNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNKnNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK`NNNNNNNNNNNNNNNNNNNNNNKuNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�K�K�K�K�K�NNNNNNNNNNNNNNNNKmNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK_NNNNNNNNNNNNNNNNNNNNNNKtNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNNKlNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK^NNNNNNNNNNNNNNNNNNNNNNKsNNNNNNNNNNNNNNNNNNNNe]�(NNNNKNNNNNNNNNNNNNNNNNNNNNKkNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK]NNNNNNNNNNNNNNNNNNNNKrKsKrKqKrNNNNNNNNNNNNNNNNNNe]�(NNNNK~NNNNNNNNNNNNNNNNNNNNNKjNNNNNNNNNNNNNNNNNNNNNNNK^K]K\K[KZK[K\K]K^NNNNNNNNNNNNNNNNNNKqKrKqKpKqNNNNNNNNNNNNNNNNNNe]�(NNNNK}NNNNNNNNNNNNNNNNNNNNNKiNNNNNNNNNNNNNNNNNNNNNNNK]K\K[KZKYKZK[K\K]NNNNNNNNNNNNNNNNNNKpKqKpKoKpNNNNNNNNNNNNNNNNNNe]�(NNNNK|NNNNNNNNNNNNNNNNNNNNKiKhKgKfKgKhKiKjKkNNNNNNNNNNNNNNNNK\K[KZKYKXKYKZK[K\NNNNNNNNNNNNNNNKlKmKnKoKpKoKnKoNNNNNNNNNNNNNNNNNNe]�(NNNNK{NNNNNNNNNNNNNNKnKmKlKkKjKiKhKgKfKeKfKgKhKiKjNNNNNNNNNNNNNNNNK[KZKYKXKWKXKYKZK[NNNNNNNNNNNNNNNKkKlKmKnKoKnKmKnNNNNNNNNNNNNNNNNNNe]�(NNK|K{KzK{K|K}K~KK�NNNNNNNNKoNNNNNKgKfKeKdKeKfKgKhKiNNNNNNNNNNNNNNNNKZKYKXKWKVKWKXKYKZNNNNNNNNNKdKeKfKgKhKiKjKkKlKmKnKmKlKmNNNNNNNNNNNNNNNNNNe]�(NNK{KzKyKzK{K|K}K~KNNNNNNNNKpNNNNNKfKeKdKcKdKeKfKgKhNNNNNNNNNNNNNNNNKYKXKWKVKUKVKWKXKYKZK[K\K]K^K_K`KaKbKcNNNNNKkKlKmKnKmKlKkKlNNNNNNNNNNNNNNNNNNe]�(NNKzKyKxKyKzK{K|K}K~NNNNNNNNKqNNNNNKeKdKcKbKcKdKeKfKgNNNNNNNNNNNNNNNNKXKWKVKUKTKUKVKWKXNNNNNNNNNNNNNNNKlKmKnKmKlKkKjKkNNNNNNNNNNNNNNNNNNe]�(NNKyKxKwNNKzK{K|K}NNNNNNNNKrNNNNNKdKcKbKaKbKcKdKeKfNNNNNNNNNNNNNNNNKWKVKUKTKSKTKUKVKWNNNNNNNNNNNNNNNNNNNNNKiNNNNNNNNNNNNNNNNNNNe]�(NNKxKwKvNNKyKzK{K|NNNNNNNNKsNNNNNKcKbKaK`KaKbKcKdKeNNNNNNNNNNNNNNNNKVKUKTKSKRKSKTKUKVNNNNNNNNNNNNNNNNNNNNNKhNNNNNNNNNNNNNNNNNNNe]�(NNKwKvKuKvKwKxKyKzK{NNNNNNNNKtNNNNNKbKaK`K_K`KaKbKcKdNNNNNNNNNNNNNNNNKUKTKSKRKQKRKSKTKUNNNNNNNNNNNNNNNNNNNNNKgNNNNNNNNNNNNNNNNNNNe]�(NNKvKuKtKuKvKwKxKyKzNNNNNNNNKuNNNNNKaK`K_K^K_K`KaKbKcNNNNNNNNNNNNNNNNNNNNKPNNNNNNNNNNNNNNNK\K]K^K_K`KaKbKcKdKeKfNNNNNNNNNNNNNNNNNNNe]�(NNKuKtKsKtKuKvKwKxKyKzK{K|K{KzKyKxKwKvNNNNNK`K_K^K]K^K_K`KaKbNNNNNNNNNNNNNNNNNNNNKONNNNNNNNNNNNNNNK[NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKrNNNNNNNNNNNNNNNNNNNNNNNK\NNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKZNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKqKpKoKnKmNNNNNNNNNNNNNNNNNNNK[NNNNNNNNNNNNNNNNNNNNNNNNNKMKLKKKJKINNNNNNNNNNNKYNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKlNNNNNNNNNNNNNNNNNNNKZNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKHNNNNNNNNNNNKXNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKkNNNNNNNNNNNNNNNNNNNKYKXKWKVKUNNNNNNNNNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNKWNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKpKoKnKmKlKkKjKiKhKgNNNNNNNNNNNNNNNNNNNNKTNNNNNNNNNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNKVNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKoKnKmKlKkKjKiKhKgKfNNNNNNNNNNNNNNNNNNNNKSNNNNNNNNNNNNNNNNNNNNNNNNNKENNNNNNNNNNKTKUKVKWKXKYKZK[K\NNNNNNNNNNNNNNNNNNNNNNe]�(NNKnKmKlKkKjKiKhKgKfKeKdKcKbKaK`K_K^K]NNNNNNNNNKSKRKQKRKSNNNNNNNNNNNNNNNNNNNNNNNNKDNNNNNNNNNNKSKTKUKVKWKXKYKZK[NNNNNNNNNNNNNNNNNNNNNNe]�(NNKoKnKmKlKkKjKiKhKgKfNNNNNNNK\NNNNNNNNNKRKQKPKQKRNNNNNNNNNNNNNNNNNNK?K>K?K@KAKBKCNNNNNNNNNNKRKSKTKUKVKWKXKYKZNNNNNNNNNNNNNNNNNNNNNNe]�(NNKpKoKnKmKlKkNNNKgNNNNNNNK[NNNNNNNKSKRKQKPKOKPKQNNNNNNNNNNNNNNNNNNK>K=K>K?K@KAKBKCKDKEKFKGKHKIKJNNKQKRKSKTKUKVKWKXKYNNNNNNNNNNNNNNNNNNNNNNe]�(NNKqKpKoKnKmKlNNNKhNNNNNNNKZNNNNNNNKRKQKPKOKNKOKPNNNNNNNNNNNNNNNNNNK=K<K=K>K?K@KANNNNNNNKKNNKPKQKRKSKTKUKVKWKXNNNNNNNNNNNNNNNNNNNNNNe]�(NNKrKqKpKoKnKmNNNKiNNNNNNNKYKXKWKVKUKTKSKRKQKPKOKNKMKNKONNNNNNNNNNNNNNNNNNK<K;K<K=K>K?K@NNNNNNNKLKMKNKOKPKQKRKSKTKUKVKWNNNNNNNNNNNNNNNNNNNNNNe]�(NNKsKrKqKpKoKnKmKlKkKjNNNNNNNNNNNNNNNKPKOKNKMKLKMKNNNNNNNNNNNNNNNNNNNK;K:K;K<K=K>K?NNNNNNNNNNKPKQKRKSKTKUKVKWKXNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKpNNNNNNNNNNNNNNNNNNNNKOKNKMKLKKKLKMNNNNNNNNNNNNNNNNNNK:K9K:K;K<K=K>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKqNNNNNNNNNNNNNNNNNNNNNNNNKJNNNNNNNNNNNNNNNNNNNNK9K8K9K:K;K<K=NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKrNNNNNNNNNNNNNNNNNNNNNNNNKINNNNNNNNNNNNNNNNNNNNK8K7K8K9K:K;K<NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKqNNNNNNNNNNNNNNNNNNNNNNNNKHNNNNNNNNNNNNNNNNNNNNK7K6K7K8K9K:K;NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKpNNNNNNNNNNNNNNNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNK6K5K6K7K8K9K:NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKlKmKnKoNNNNNNNNNNNNNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKkNNNNNNNNNNNNNNNNNNNNNNNNNNNKENNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKjNNNNNNNNNNNNNNNNNNNNNNNNNKBKCKDNNNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKiNNNNNNNNNNNNNNNNNNNNNNNNNKANNNNNNNNNNNNNNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKhNNNNNNNNNNNNNNNNNNNNNNNNNK@NNNNNNNNNNNNNNNNNK*K+K,K-K.K/K0NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKgNNNNNNNNNNNNNNNNNNNNNKCKBKAK@K?K>K=K<NNNNNNNNNNNNNNK)NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKgKfKeKdKcKbKaNNNNNNNNNNNNNNNNKBKAK@K?K>K=K<K;K:K9K8K7K6NNNNNNNNNK(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKfKeKdKcKbKaK`NNNNNNNNNNNNNNNNKCKBKAK@K?K>K=K<NNNNK5NNNNNNNNNK'NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKeKdKcKbKaK`K_NNNNNNNNNNNNNNNNKDKCNNNK?K>K=NNNNK4NNNNNNNNNK&NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKdKcKbKaK`K_K^NNNNNNNNNNNNNNNNKEKDNNNK@K?K>NNNNK3NNNNNNNNK&K%K$K#K"K!K KNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKcKbKaK`K_K^K]NNNNNNNNNNNNNNNNKFKENNNKAK@K?NNNNK2NNNNNNNNK%K$K#K"K!K KKNNNNNNNNNNNNNNNNNKKK
K	KKKKKKNNNNNNNNNNNNNNNNNNNe]�(NNKbKaK`K_K^K]K\NNNNNNNNKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@NNNNK1NNNNNNNNK$K#K"K!K KKKNNNNNNNNNNNNNNNNNKK
K	KKKKKKKNNNNNNNNNNNNNNNNNNNe]�(NNKcKbNNK]K\K[NNNNNNNNKPNNNNNNNKHKGKFKEKDKCKBKANNNNK0NNNNNNNNK#K"K!K KKKKKKKKKKKKKKKNNNNNNK
K	KKKKKKKKNNNNNNNNNNNNNNNNNNNe]�(NNKbKaNNK\K[KZKYKXKWKVKUKTKSKRKQNNNNNNNNNNNNNNNNNNNK/NNNNNNNNK$K#K"K!K KKKNNNNNNNNNNKKKKKKK
K	KKKKKKKKKNNNNNNNNNNNNNNNNNNNe]�(NNKaK`K_K^K]K\K[NNNNNNNNNNNNNNNNNNNNNNNNNNNNK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKNNNNNNNNNNNNNNNNNKKKKKKKKK KNNNNNNNNNNNNNNNNNNNe]�(NNKbKaK`K_K^K]K\NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK#K"K!K KNNNNNNNNNNNNNNNNNK	KKKKKKKKKNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK$K#K"K!K NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK%K$K#K"K!NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeehA�1A: Sacked Tower�j  }�(Kj�  )��}�(j�  KJj�  j�  j�  �Features.Features��Chest���)��}�(h^jw~  hDhEhV]�hj�}  hAjz~  ubj  K�ID�Khj�}  hAjz~  ubKj�  )��}�(j�  KGj�  j�  j�  j{~  )��}�(h^j�~  hDhEhV]�hj�}  hAjz~  ubj  Kj~  Khj�}  hAjz~  ubKj�  )��}�(j�  KNj�  j�  j�  j  j  K	j~  KhhChA�Item�ubKj�  )��}�(j�  Kj�  j�  j�  j{~  )��}�(h^j�~  hDhEhV]�hj�}  hAjz~  ubj  Kj~  Khj�}  hAjz~  ubKj�  )��}�(j�  Kj�  j�  j�  j{~  )��}�(h^j�~  hDhEhV]�hj�}  hAjz~  ubj  Kj~  Khj�}  hAjz~  ubKj�  )��}�(j�  K
j�  j�  j�  j  )��}�(h^Nh>h<hD]�(K�K�KehG�h<��coins�Kh�$�hA�
Gold Coins�ubj  Kj~  Khji  hA�Health�ubK#j�  )��}�(j�  K6j�  j�  j�  jy~  �Brush���)��}�(h^j�~  hD]�(KKnKehj�}  hAj�~  ubj  K#j~  K#hj�}  hAj�~  ubK$j�  )��}�(j�  K7j�  j�  j�  j�~  )��}�(h^j�~  hDj�~  hj�}  hAj�~  ubj  K#j~  K$hj�}  hAj�~  ubK&j�  )��}�(j�  K8j�  j�  j�  h�j  K(j~  K&hji  hAj�~  ubK'j�  )��}�(j�  KNj�  j�  j�  j{~  )��}�(h^j�~  hDhEhV]�hj�}  hAjz~  ubj  K(j~  K'hj�}  hAjz~  ubK*j�  )��}�(j�  KNj�  j�  j�  j{~  )��}�(h^j�~  hDhEhV]�hj�}  hAjz~  ubj  K)j~  K*hj�}  hAjz~  ubK,j�  )��}�(j�  K9j�  j�  j�  j{~  )��}�(h^j�~  hDhEhV]�hj�}  hAjz~  ubj  K+j~  K,hj�}  hAjz~  ubK.j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(�
stealthVal�K hK �isAfraid��hKhKh]�hNh1�h-Kh.K �	cowardice�G?�      �
dropChance�K(j�  Kh/�h0NhKd�
alliesList�]�(j�~  j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�      j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�~  j�~  j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�      j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�~  j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�      j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�~  j�~  j�~  j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�      j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�~  j�~  j�~  j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�������j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�~  j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G        j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�~  j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�������j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�~  j�~  j�~  eh3�h6j�|  )��}�(h<�h-K h=Kh_Kh>h?h@�hKhAj�|  hB�hKhhChDhEhF�hG�hHK ubhIKhJ�hLK hMhj)��}�(h<�h-Kh=Kh>hRh@�hKhAhihB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUK
hV]�j�  K �hearingDist�KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  ��lastPlayerMap�NhA�Goblin Lancer�h^j�~  �necklace�N�accuracy�K hD]�(K�KKe�lastPlayerLoc�N�	sightDist�K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  KKj~  KOhj�}  hA�Enemy�ubj�~  eh3�h6j  )��}�(h<�h-K h=Kh_Kh>hvh@�hKhAj  hB�hKhhChDhEhF�hG�hHK ubhIKhJ�hLK hMh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hej�|  )��}�(h=K7hKh>hehDhEhF�hG�h<�h_K2hhChA�Iron Breastplate�ubhj�}  j�  �j�~  NhA�Goblin Stonewall�h^j�~  j�~  Nj�~  K hDj�~  j�~  Nj�~  Kh_K h]hn)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAhqububj  KKj~  KNhj�}  hAj�~  ubj�~  j�~  eh3�h6j�|  )��}�(h<�h-K h=Kh_Kh>h?h@�hKhAj�|  hB�hKhhChDhEhF�hG�hHK ubhIKhJ�hLK hMhj)��}�(h<�h-Kh=Kh>hRh@�hKhAhihB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj�~  h^j�~  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  KNj~  KRhj�}  hAj�~  ubeh3�h6h�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhIKhJ�hLK hMh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKub�optionalTargets�]�j�~  j�~  ��ahS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhA�Goblin Thief�h^j�~  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  KGj~  K[hj�}  hAj�~  ubeh3�h6h�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhIKhJ�hLK hMh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubj  ]�j  ahS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj   h^j�~  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  KEj~  KKhj�}  hAj�~  ubj�~  j�~  eh3�h6h�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhIKhJ�hLK hMh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubj  ]�j  ahS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj   h^j�~  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  KEj~  KWhj�}  hAj�~  ubj�~  eh3�h6h�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhIKhJ�hLK hMh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubj  ]�j  ahS�j�  K hUKhV]�hj)��}�(h^Nh<�h-Kh=Kh>hRh@�hKhAhihB�hKhhChDhEhF�hG�hKhHKubaj�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj   h^j�~  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  KEj~  KPhj�}  hAj�~  ubeh3�h6h�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhIKhJ�hLK hMh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubj  ]�j  ahS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj   h^j�~  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  KBj~  K.hj�}  hAj�~  ubK/j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G        j�~  K(j�  Kh/�h0NhKdj�~  ]�jQ  ah3�h6j  )��}�(h<�h-K h=Kh_Kh>hvh@�hKhAj  hB�hKhhChDhEhF�hG�hHK ubhIKhJ�hLK hMh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hej�|  )��}�(h=K7hKh>hehDhEhF�hG�h<�h_K2hhChAj  ubhj�}  j�  �j�~  NhAj  h^jQ  j�~  Nj�~  K hDj�~  j�~  Nj�~  Kh_K h]hn)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAhqububj  K,j~  K/hj�}  hAj�~  ubK0j�  )��}�(j�  Kj�  j�  j�  j{~  )��}�(h^ja  hD]�(KQKOKehV]�(j
  )��}�(�
arrowCount�Kh>h<hDhEhG�h<�h�i�hA�Bundle of Arrows�ubj  )��}�(h<�h-K h=Kh_Kh>hvh@�hKhAj  hB�hKhhChDhEhF�hG�hHK ubhZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ubj  )��}�(h>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubehj�}  hAjz~  ubj  K,j~  K0hj�}  hAjz~  ubK1j�  )��}�(j�  K
j�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G        j�~  K(j�  Kh/�h0NhKdj�~  ]�(jQ  jr  j�  )��}�(j�  K
j�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G        j�~  K(j�  Kh/�h0NhKdj�~  ]�(jQ  jr  jx  eh3�h6NhIKhJ�hLK hMhO)��}�(h<�h-Kh=Kh>hRh@�hKhAhNhB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhA�Goblin Berserker�h^jx  j�~  Nj�~  K hDj�~  j�~  Nj�~  Kh_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  K0j~  K:hj�}  hAj�~  ubeh3�h6NhIKhJ�hLK hMhO)��}�(h<�h-Kh=Kh>hRh@�hKhAhNhB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUK
hV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj�  h^jr  j�~  Nj�~  K hDj�~  j�~  Nj�~  Kh_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  K,j~  K1hj�}  hAj�~  ubK3j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?��Q�j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�  j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G        j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�  j�  eh3�h6j  )��}�(h<�h-K h=Kh_Kh>hvh@�hKhAj  hB�hKhhChDhEhF�hG�hHK ubhIKhJ�hLK hMh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hej�|  )��}�(h=K7hKh>hehDhEhF�hG�h<�h_K2hhChAj  ubhj�}  j�  �j�~  NhAj  h^j�  j�~  Nj�~  K hDj�~  j�~  Nj�~  Kh_K h]hn)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAhqububj  K1j~  K=hj�}  hAj�~  ubj�  )��}�(j�  K!j�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?��Q�j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�  j�  j�  eh3�h6NhIKhJ�hLK hMhs)��}�(h<�h-Kh=Kh>hvh@�hKhAhrhB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhA�Goblin Grunt�h^j�  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  K2j~  K>hj�}  hAj�~  ubeh3�h6NhIKhJ�hLK hMhs)��}�(h<�h-Kh=Kh>hvh@�hKhAhrhB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj�  h^j�  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  K-j~  K3hj�}  hAj�~  ubK4j�  )��}�(j�  K2j�  j�  j�  h�j  K-j~  K4hhChAj�~  ubK8j�  )��}�(j�  Kj�  j�  j�  h�)��}�(h^j�  h<�h�Kh>h<hK hAh�h�KhKhh�hDhEj   KhG�j  j  ubj  K/j~  K8hji  hAj�~  ubK9j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�      j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?��Q�j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�  j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G        j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�  j�  eh3�h6j  )��}�(h<�h-K h=Kh_Kh>hvh@�hKhAj  hB�hKhhChDhEhF�hG�hHK ubhIKhJ�hLK hMh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hej�|  )��}�(h=K7hKh>hehDhEhF�hG�h<�h_K2hhChAj  ubhj�}  j�  �j�~  NhAj  h^j�  j�~  Nj�~  K hDj�~  j�~  Nj�~  Kh_K h]hn)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAhqububj  K9j~  K@hj�}  hAj�~  ubj�  j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�      j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�  j�  j�  j�  eh3�h6h�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhIKhJ�hLK hMh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubj  ]�j  ahS�j�  K hUK	hV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj   h^j�  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  K>j~  KBhj�}  hAj�~  ubeh3�h6NhIKhJ�hLK hMhs)��}�(h<�h-Kh=Kh>hvh@�hKhAhrhB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj�  h^j�  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  K9j~  K?hj�}  hAj�~  ubj�  j�  j�  eh3�h6h�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhIKhJ�hLK hMh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubj  ]�j  ahS�j�  K hUKhV]�hb)��}�(h=KhKh>heh^NhDhEhF�hG�h<�h_KhhChAhfubaj�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj   h^j�  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  K?j~  K9hj�}  hAj�~  ubK:jx  K<j�  )��}�(j�  Kj�  j�  j�  j�  j  K1j~  K<hhChAj�~  ubK=j�  K>j�  K?j�  K@j�  KBj�  KCj�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�      j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�  j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?��Q�j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�  j�  j�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�      j�~  K(j�  Kh/�h0NhKdj�~  ]�(j�  j�  j�  eh3�h6NhIKhJ�hLKhMh�)��}�(h<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhA�Goblin Archer�h^j�  j�~  Nj�~  K hDj�~  j�~  Nj�~  K
h_K h]h)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAh�ububj  K?j~  KLhj�}  hAj�~  ubeh3�h6NhIKhJ�hLK hMhs)��}�(h<�h-Kh=Kh>hvh@�hKhAhrhB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj�  h^j�  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  K=j~  KHhj�}  hAj�~  ubj�  eh3�h6NhIKhJ�hLKhMh�)��}�(h<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj�  h^j�  j�~  Nj�~  K hDj�~  j�~  Nj�~  K
h_K h]h)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAh�ububj  K:j~  KChj�}  hAj�~  ubKDj�  )��}�(j�  KLj�  j�  j�  j{~  )��}�(h^j1�  hDhEhV]�hj�}  hAjz~  ubj  K;j~  KDhj�}  hAjz~  ubKEj�  )��}�(j�  K9j�  j�  j�  �Features.Stairs��StairUp���)��}�(j�  K9j�  j�  h^j6�  j�  Nj  K<j~  J�����moveCost�KhA�Stairs�ubj  K<j~  KEhj�}  hA�	Stairs Up�ubKFj�  KGj�  )��}�(j�  K5j�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�      j�~  K(j�  Kh/�h0NhKdj�~  ]�j@�  ah3�h6h�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhIKhJ�hLK hMh�)��}�(h<�h-Kh=Kh>hvh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubj  ]�j  ahS�j�  K hUK
hV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK\K[KZKYNNNNNNNNNNNNNNNNNKGKHKIKJKKKLNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK[KZKYKXNNNNNNNNNNNNNNNNNKFKGKHKIKJKKNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�KNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK\K[KZKYKXKWNNNNNNNNNNNNNNNNNKEKFKGKHKIKJNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�KK~K}K|K{KzKyKxKwKvKuNNNNNNNNNNNNNNNNNNNKaK`K_K^K]K\K[KZKYKXKWKVNNNNNNNNNNNNNNNNNKDKEKFKGKHKIKJKKKLNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�KNNNNNNNNKtNNNNNNNNNNNNNNNNNNNKbNNNNNKZKYKXKWKVKUNNNNNNNNNNNNNNNNNKCKDKEKFKGKHKIKJKKNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNKsNNNNNNNNNNNNNNNNNNNKcNNNNNKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJNNNNNNNKBKCKDKEKFKGKHKIKJNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNKrNNNNKmKlKkKjKkKlNNNNNNNNNKdNNNNNKZNNNNNNNNNNNNNNKIKHKGKFKEKDKCKBKAKBKCKDKEKFKGKHKINNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNKqKpKoKnKmKlKkKjKiKjKkKlKmKlKkKjKiKhKgKfKeNNNNNK[NNNNNNNNNNNNNNNNNNNNNNK@KAKBKCKDKEKFKGKHNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNKkKjKiKhNNNNNNNNNNNNNNNNNKZNNNNNNNNNNNNNNNNNNNNNNK?NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNKjKiKhKgNNNNNNNNNNNNNNNNNKYNNNNNNNNNNNNNNNNNNNNNNK>NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK�K�K�K�K�K�K�NNNNNNNNNNNNNKiKhKgKfKgKhNNNNNNNNNNNNNNNKXNNNNNNNNNNNNNNNNNNNNNNK=NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNKhKgKfKeKfKgNNNNNNNNNNNNNNNKWNNNNNNNNNNNNNNNNNNNNNNK<NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNKgKfKeKdKeKfNNNNNNNNNNNNNNNKVNNNNNNNNNNNNNNNNNNNNNNK;NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNKfKeKdKcKdKeNNNNNNNNNNNNNNNKUNNNNNNNNNNNNNNNNNNNNNNK:NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNKbNNNNNNNNNNNNNNNNNKTKSKRKQKPKOKNNNNNNNNNNNNNNNNNK9NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNKaNNNNNNNNNNNNNNNNNNNNNNNKMNNNNNNNNNNNNNNNNK8NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNK`NNNNNNNNNNNNNNNNNNNNNNNKLNNNNNNNNNNNNNNNNK7NNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNK_K^NNNNNNNNNNNNNNNNNNNNNNKKNNNNNNNNNNNNNNNNK6K5K4NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK�NNNNNNNNNNNNNNNNNNNNNK]NNNNNNNNNNNNNNNNNNNNNNKJNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�K�K�K�NNNNNNNNNNNNNNNNNNNNNK\NNNNNNNNNNNNNNNNNNNNNNKINNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNKaK`K_K^K]K\K[KZKYKXNNNNNNNNNNNNNNNNNNNKHNNNNNNNNNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKONNNNNNNNNNNKGNNNNNNNNNNNNNNNNNNK0NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNKaK`K_K^K]K\K[KZKYKXNNNNNNNKNNNNNNNNNNNNKFNNNNNNNNNNNNNNNNNNK/NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNKbKaK`NNNNK[KZKYNNNNNNNKMNNNNNNNNNNNKENNNNNNNNNNNNNNNNK0K/K.K-K,K-K.K/K0K1NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNNNNNNNKcKbKaNNNNK\K[KZNNNNNNNKLNNNNNNNNKCKBKCKDKEKFKGKHKGNNNNNNNNK2K1K0K/K.K-K,K+K,K-K.K/K0NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�KNNNNNNNNKjKiKhKgKfKeKdKcKbNNNNK]K\K[NNNNNNNKKNNNNNNNNKBKAKBKCKDKEKFKGKFNNNNNNNNK3NNK.K-K,K+K*K+K,K-K.K/NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�KK~NNNNNNNNKkNNNNNKeKdKcNNNNK^K]K\NNNNNNNKJKIKHKGKFKEKDKCKBKAK@KAKBKCKDKEKFKENNNNNNNNK4NNK-K,K+K*K)K*K+K,K-K.NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�KK~K}NNNNNNNNKlNNNNNKfKeKdKcKbKaK`K_K^K]NNNNNNNNNNNNNNNNK@K?K@KAKBKCKDKEKDNNNNNNNNK5NNNNK*K)K(K)K*K+K,K-NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK}K|NNNNNNNNKmNNNNNKgKfKeKdKcKbKaK`K_K^NNNNNNNNNNNNNNNNK?K>K?K@KAKBKCKDKCNNNNNNNNK6NNNNK)K(K'K(K)K*K+K,NNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK|K{NNNNNNNNKnNNNNNNKgNNNNNNNNNNNNNNNNNNNNNNNNK>K=K>K?K@KAKBKCKBNNNNNNNNK7NNNNNNK&NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNK{KzNNNNNNNNKoNNNNNNKhNNNNNNNNNNNNNNNNNNNNNNNNK=K<K=K>K?K@KAKBKAK@K?K>K=K<K;K:K9K8NNNNNNK%NNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNNNKzKyKxKwKvKuKtKsKrKqKpNNNNNNKiNNNNNNNNNNNNNNNNNNNNNNNNNK;NNNNNNNNNNNNNNNNNNNNNNK$K#K"K!K NNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK{NNNNNNNNNNNNNNNNKjNNNNNNNNNNNNNNNNNNNNNNNNNK:NNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK|NNNNNNNNNNNNNNNNKkNNNNNNNNNNNNNNNNNNNNNNNNNK9K8K7K6K5NNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK}NNNNNNNNNNNNNNNNKlNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�K�K�K�KK~NNNNNNNNNNNNNNNNKmNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNNKnNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNNKoNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNNKpNNNNNNNNNNNNNNNNNNNNNNNK2K1K0K/K.K/K0K1K0NNNNNNNNNNNNNNNNNNKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNNKqNNNNNNNNNNNNNNNNNNNNNNNK1K0K/K.K-K.K/K0K/NNNNNNNNNNNNNNNNNNKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNKsKrKsKtKuKvKwKxKyNNNNNNNNNNNNNNNNK0K/K.K-K,K-K.K/K.NNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNKzKyKxKwKvKuKtKsKtKuKvKwKxKyKzNNNNNNNNNNNNNNNNK/K.K-K,K+K,K-K.K-NNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK{NNNNNKuKtKuKvKwKxKyKzK{NNNNNNNNNNNNNNNNK.K-K,K+K*K+K,K-K,NNNNNNNNNK KKKKKKKKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK|NNNNNKvKuKvKwKxKyKzK{K|NNNNNNNNNNNNNNNNK-K,K+K*K)K*K+K,K+K*K)K(K'K&K%K$K#K"K!NNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK}NNNNNKwKvKwKvKwKxKyKzK{NNNNNNNNNNNNNNNNK,K+K*K)K(K)K*K+K,NNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNK�K�K�K�NNNNNNNNK~NNNNNKxKwKvKuKvKwKxKyKzNNNNNNNNNNNNNNNNK+K*K)K(K'K(K)K*K+NNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�NNK�K�K�K�NNNNNNNNKNNNNNKwKvKuKtKuKvKwKxKyNNNNNNNNNNNNNNNNK*K)K(K'K&K'K(K)K*NNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK�NNNNNKvKuKtKsKtKuKvKwKxNNNNNNNNNNNNNNNNK)K(K'K&K%K&K'K(K)NNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�NNNNNNNNK�NNNNNKuKtKsKrKsKtKuKvKwNNNNNNNNNNNNNNNNNNNNK$NNNNNNNNNNNNNNNKKKKKK	K
KKKKNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�K�NNNNNKtKsKrKqKrKsKtKuKvNNNNNNNNNNNNNNNNNNNNK#NNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�NNNNNNNNNNNNNNNNNNNNNNNKpNNNNNNNNNNNNNNNNNNNNNNNNNK"NNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNK�K�K�K�K�NNNNNNNNNNNNNNNNNNNKoNNNNNNNNNNNNNNNNNNNNNNNNNK!K KKKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNK�NNNNNNNNNNNNNNNNNNNKnNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNK NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNKNNNNNNNNNNNNNNNNNNNKmKlKkKjKiNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�KK~K}K|K{NNNNNNNNNNNNNNNNNNNNKhNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�KK~K}K|K{KzNNNNNNNNNNNNNNNNNNNNKgNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNKKKKKKKK	K
NNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�KK~K}K|K{KzKyKxKwKvKuKtKsKrKqNNNNNNNNNKgKfKeKfKgNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNKKKKKKK	K
KNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�KK~K}K|K{KzNNNNNNNKpNNNNNNNNNKfKeKdKeKfNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNKKKKKK	K
KKNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�KNNNK{NNNNNNNKoNNNNNNNKgKfKeKdKcKdKeNNNNNNNNNNNNNNNNNNKKKKKKKKKKKKKKKNNKKKKK	K
KKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�NNNK|NNNNNNNKnNNNNNNNKfKeKdKcKbKcKdNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNKNNKKKK	K
KKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�NNNK}NNNNNNNKmKlKkKjKiKhKgKfKeKdKcKbKaKbKcNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNKKK
K	KK	K
KKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNK�K�K�K�K�K�K�K�KK~NNNNNNNNNNNNNNNKdKcKbKaK`KaKbNNNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNK
K	K
KKKKKKNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNNNKcKbKaK`K_K`KaNNNNNNNNNNNNNNNNNNK KKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNK^NNNNNNNNNNNNNNNNNNNNK!K KKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNK]NNNNNNNNNNNNNNNNNNNNK"K!K KKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNK\NNNNNNNNNNNNNNNNNNNNK#K"K!K KKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK�NNNNNNNNNNNNNNNNNNNNNNNNK[NNNNNNNNNNNNNNNNNNNNK$K#K"K!K KKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNK�K�K�K�NNNNNNNNNNNNNNNNNNNNNNNNKZNNNNNNNNNNNNNNNNNNNNNK$NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNKYNNNNNNNNNNNNNNNNNNNNNK%NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNK~NNNNNNNNNNNNNNNNNNNNNNNNNKVKWKXNNNNNNNNNNNNNNNNNNNNNK&NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNK}NNNNNNNNNNNNNNNNNNNNNNNNNKUNNNNNNNNNNNNNNNNNNNNNNNK'NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNK|NNNNNNNNNNNNNNNNNNNNNNNNNKTNNNNNNNNNNNNNNNNNK.K-K,K+K*K)K(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNK{NNNNNNNNNNNNNNNNNNNNNKWKVKUKTKSKRKQKPNNNNNNNNNNNNNNK/NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK{KzKyKxKwKvKuNNNNNNNNNNNNNNNNKVKUKTKSKRKQKPKOKNKMKLKKKJNNNNNNNNNK0NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKzKyKxKwKvKuKtNNNNNNNNNNNNNNNNKWKVKUKTKSKRKQKPNNNNKINNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKyKxKwKvKuKtKsNNNNNNNNNNNNNNNNKXKWNNNKSKRKQNNNNKHNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKxKwKvKuKtKsKrNNNNNNNNNNNNNNNNKYKXNNNKTKSKRNNNNKGNNNNNNNNK4K3K4K5K6K7K8K9NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKwKvKuKtKsKrKqNNNNNNNNNNNNNNNNKZKYNNNKUKTKSNNNNKFNNNNNNNNK5K4K5K6K7K8K9K:NNNNNNNNNNNNNNNNNKRKSKTKUKVKWKXKYKZK[NNNNNNNNNNNNNNNNNNNe]�(NNKvKuKtKsKrKqKpNNNNNNNNKcKbKaK`K_K^K]K\K[KZKYKXKWKVKUKTNNNNKENNNNNNNNK6K5K6K7K8K9K:K;NNNNNNNNNNNNNNNNNKQKRKSKTKUKVKWKXKYKZNNNNNNNNNNNNNNNNNNNe]�(NNKwKvNNKqKpKoNNNNNNNNKdNNNNNNNK\K[KZKYKXKWKVKUNNNNKDNNNNNNNNK7K6K7K8K9K:K;K<K=K>K?K@KAKBKCKDKEKFKGNNNNNNKPKQKRKSKTKUKVKWKXKYNNNNNNNNNNNNNNNNNNNe]�(NNKvKuNNKpKoKnKmKlKkKjKiKhKgKfKeNNNNNNNNNNNNNNNNNNNKCNNNNNNNNK8K7K8K9K:K;K<K=NNNNNNNNNNKHKIKJKKKLKMKNKOKPKQKRKSKTKUKVKWKXNNNNNNNNNNNNNNNNNNNe]�(NNKuKtKsKrKqKpKoNNNNNNNNNNNNNNNNNNNNNNNNNNNNKBKAK@K?K>K=K<K;K:K9K8K9K:K;K<K=K>NNNNNNNNNNNNNNNNNKPKQKRKSKTKUKVKWKXKYNNNNNNNNNNNNNNNNNNNe]�(NNKvKuKtKsKrKqKpNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK;K<K=K>K?NNNNNNNNNNNNNNNNNKQKRKSKTKUKVKWKXKYKZNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK<K=K>K?K@NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK=K>K?K@KANNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeehAj   h^j@�  j�~  Nj�~  K hDj�~  j�~  ]�(K6KFej�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  Kj~  KGhj�}  hAj�~  ubKHj�  KKj�~  KLj�  KMj�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�      j�~  K(j�  Kh/�h0NhKdj�~  ]�j��  ah3�h6NhIKhJ�hLKhMh�)��}�(h<�h-Kh=Kh>hRh@�hKhAh�hB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj�  h^j��  j�~  Nj�~  K hDj�~  j�~  Nj�~  K
h_K h]h)��}�(h=KhKh>h]hDhEhF�hG�h<�h_KhhChAh�ububj  KJj~  KMhj�}  hAj�~  ubKNj�~  KOj�~  KPj�~  KQj�  )��}�(j�  Kj�  j�  j�  j{~  )��}�(h^jŀ  hDje  hV]�(j  )��}�(h>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubh�)��}�(hKh>h�hDhEhG�h<�hh�h�hhAh�ubj�|  )��}�(h<�h-Kh=Kh>hRh@�hKhAj�|  hB�hKhhChDhEhF�hG�hKhHKubj  )��}�(h>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubehj�}  hAjz~  ubj  KMj~  KQhj�}  hAjz~  ubKRj�~  KSj�  )��}�(j�  Kj�  j�  j�  j{~  )��}�(h^jҀ  hDje  hV]�(h�)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAh�ubhZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ubjf  )��}�(h>h<hDhEhG�h<�hji  jj  KhAjk  ubj  )��}�(h>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubehj�}  hAjz~  ubj  KNj~  KShj�}  hAjz~  ubKTj�  )��}�(j�  Kj�  j�  j�  j~  )��}�(j�~  K hK j�~  �hKhKh]�hNh1�h-Kh.K j�~  G?�������j�~  K(j�  Kh/�h0NhKdj�~  ]�j߀  ah3�h6j�|  )��}�(h<�h-K h=Kh_Kh>h?h@�hKhAj�|  hB�hKhhChDhEhF�hG�hHK ubhIKhJ�hLK hMhj)��}�(h<�h-Kh=Kh>hRh@�hKhAhihB�hKhhChDhEhF�hG�hKhHKubhS�j�  K hUKhV]�j�  K j�~  KhTKj�  ]�hehb)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAhfubhj�}  j�  �j�~  NhAj�~  h^j߀  j�~  Nj�~  K hDj�~  j�~  Nj�~  K	h_K h]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ububj  KOj~  KThj�}  hAj�~  ubKVj�  )��}�(j�  KLj�  j�  j�  j{~  )��}�(h^j�  hDje  hV]�(hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ubj�|  )��}�(h<�h-Kh=Kh>hRh@�hKhAj�|  hB�hKhhChDhEhF�hG�hKhHKubh�)��}�(h<�h�Kh>h<hK hAh�h�KhKhh�hDhEj   KhG�j  j  ubj  )��}�(h>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubehj�}  hAjz~  ubj  KOj~  KVhj�}  hAjz~  ubKWj�~  KXj�  )��}�(j�  Kj�  j�  j�  j�~  )��}�(h^j��  hDj�~  hj�}  hAj�~  ubj  KPj~  KXhj�}  hAj�~  ubKYj�  )��}�(j�  Kj�  j�  j�  j�~  )��}�(h^j �  hDj�~  hj�}  hAj�~  ubj  KPj~  KYhj�}  hAj�~  ubKZj�  )��}�(j�  Kj�  j�  j�  j�~  )��}�(h^j�  hDj�~  hj�}  hAj�~  ubj  KPj~  KZhj�}  hAj�~  ubK[j�~  K]j�  )��}�(j�  Kj�  j�  j�  j�~  )��}�(h^j�  hDj�~  hj�}  hAj�~  ubj  KQj~  K]hj�}  hAj�~  ubKbj�  )��}�(j�  Kj�  j�  j�  j�~  )��}�(h^j�  hDj�~  hj�}  hAj�~  ubj  KRj~  Kbhj�}  hAj�~  ubKcj�  )��}�(j�  Kj�  j�  j�  j�~  )��}�(h^j�  hDj�~  hj�}  hAj�~  ubj  KRj~  Kchj�}  hAj�~  ubKdj�  )��}�(j�  Kj�  j�  j�  j�~  )��}�(h^j�  hDj�~  hj�}  hAj�~  ubj  KRj~  Kdhj�}  hAj�~  ubKfj�  )��}�(j�  KPj�  j�  j�  j�|  )��}�(h^j�  )��}�(j�  KFj�  j�  j�  j�  j  KRj~  K�hhChAj�|  ubh<�h-K h=Kh_Kh>h?h@�hKhAj�|  hB�hKhhChDhEhF�hG�hHK ubj  KRj~  KfhhChAj�~  ubKhj�  )��}�(j�  KOj�  j�  j�  j8�  �	StairDown���)��}�(j�  KOj�  j�  h^j�  j�  Nj  KSj~  J����hAj>�  j=�  Kubj  KSj~  Khhj�}  hA�Stairs Down�ubKij�  )��}�(j�  Kj�  j�  j�  j?  j  KTj~  KihhChAj�~  ubKjj�  )��}�(j�  K6j�  j�  j�  h[j  K3j~  KjhhChAh`ubKkj�  )��}�(j�  K6j�  j�  j�  hkj  K3j~  KkhhChAhiubKlj�  )��}�(j�  K6j�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  K3j~  Klhj�~  hAj�~  ubKmj�  )��}�(j�  K6j�  j�  j�  h[j  K3j~  KmhhChAh`ubKnj�  )��}�(j�  K6j�  j�  j�  hcj  K3j~  KnhhChAhfubKoj�  )��}�(j�  K6j�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  K3j~  Kohj�~  hAj�~  ubKpj�  )��}�(j�  K6j�  j�  j�  hkj  K3j~  KphhChAhiubKqj�  )��}�(j�  K6j�  j�  j�  hgj  K3j~  KqhhChAhfubKrj�  )��}�(j�  K6j�  j�  j�  j
  )��}�(ji  Kh>h<h^NhDhEhG�h<�hjj  hAjk  ubj  K3j~  Krhjj  hAjk  ubKsj�  )��}�(j�  K6j�  j�  j�  hkj  K3j~  KshhChAhiubKtj�  )��}�(j�  K6j�  j�  j�  hwj  K3j~  KthhChAhfubKuj�  )��}�(j�  K6j�  j�  j�  h{j  K3j~  KuhhChAh}ubKvj�  )��}�(j�  K6j�  j�  j�  hoj  K2j~  KvhhChAhqubKwj�  )��}�(j�  K6j�  j�  j�  htj  K2j~  KwhhChAhrubKxj�  )��}�(j�  K6j�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  K2j~  Kxhj�~  hAj�~  ubKyj�  )��}�(j�  K4j�  j�  j�  h�j  K!j~  KyhhChAhqubKzj�  )��}�(j�  K4j�  j�  j�  h�j  K!j~  KzhhChAhrubK{j�  )��}�(j�  K4j�  j�  j�  j
  )��}�(ji  Kh>h<h^NhDhEhG�h<�hjj  hAjk  ubj  K!j~  K{hjj  hAjk  ubK|j�  )��}�(j�  K4j�  j�  j�  h�j  Kj~  K|hhChAh�ubK}j�  )��}�(j�  K4j�  j�  j�  h�j  Kj~  K}hhChAh�ubK~j�  )��}�(j�  K4j�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K~hj�~  hAj�~  ubKj�  )��}�(j�  K5j�  j�  j�  h�j  Kj~  KhhChAh�ubK�j�  )��}�(j�  K5j�  j�  j�  h�j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  K5j�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  K!j�  j�  j�  h�j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  K!j�  j�  j�  h�j  Kj~  K�hhChAhrubK�j�  )��}�(j�  K!j�  j�  j�  h�j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  K!j�  j�  j�  h�j  Kj~  K�hhChAhfubK�j�  )��}�(j�  K!j�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  K j�  j�  j�  h�j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  K j�  j�  j�  h�j  Kj~  K�hhChAhNubK�j�  )��}�(j�  K j�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAhiubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hh�hAh�ubK�j�  )��}�(j�  K
j�  j�  j�  h�j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  K
j�  j�  j�  h�j  Kj~  K�hhChAhNubK�j�  )��}�(j�  K
j�  j�  j�  h�j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  K
j�  j�  j�  h�j  Kj~  K�hhChAhfubK�j�  )��}�(j�  K
j�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAhiubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAhfubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAh}ubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  K	j�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAhiubK�j�  )��}�(j�  K	j�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAhqubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  K	j�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAhqubK�j�  )��}�(j�  K	j�  j�  j�  h�j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  K	j�  j�  j�  j
  )��}�(ji  Kh>h<h^NhDhEhG�h<�hjj  hAjk  ubj  Kj~  K�hjj  hAjk  ubK�j�  )��}�(j�  Kj�  j�  j�  h�j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  Kj�  j�  j�  h�j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  Kj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  Kj�  j�  j�  h�j  K	j~  K�hhChAh`ubK�j�  )��}�(j�  Kj�  j�  j�  h�j  K	j~  K�hhChAhNubK�j�  )��}�(j�  Kj�  j�  j�  h�j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  Kj�  j�  j�  h�j  Kj~  K�hhChAhiubK�j�  )��}�(j�  Kj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  K/j�  j�  j�  h�j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  K/j�  j�  j�  h�j  Kj~  K�hhChAhrubK�j�  )��}�(j�  K3j�  j�  j�  h�j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  K3j�  j�  j�  h�j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  K3j�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  KGj�  j�  j�  h�j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  KGj�  j�  j�  h�j  Kj~  K�hhChAhrubK�j�  )��}�(j�  KHj�  j�  j�  j  j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  KHj�  j�  j�  j
  j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  KKj�  j�  j�  j  j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  KKj�  j�  j�  j  j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  KKj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  KOj�  j�  j�  j  j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  KOj�  j�  j�  j  j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  KOj�  j�  j�  j
  )��}�(ji  Kh>h<h^NhDhEhG�h<�hjj  hAjk  ubj  Kj~  K�hjj  hAjk  ubK�j�  )��}�(j�  KOj�  j�  j�  j  j  K	j~  K�hhChAj  ubK�j�  )��}�(j�  KOj�  j�  j�  j  j  K	j~  K�hhChAhfubK�j�  )��}�(j�  KOj�  j�  j�  j!  j  K	j~  K�hhChAh�ubK�j�  )��}�(j�  KGj�  j�  j�  j#  j  K
j~  K�hhChAh`ubK�j�  )��}�(j�  KGj�  j�  j�  j-  j  K
j~  K�hhChAhNubK�j�  )��}�(j�  KGj�  j�  j�  j%  j  Kj~  K�hhChAhqubK�j�  )��}�(j�  KGj�  j�  j�  j+  j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  KGj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  KGj�  j�  j�  j'  j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  KGj�  j�  j�  j)  j  Kj~  K�hhChAhrubK�j�  )��}�(j�  KGj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  KHj�  j�  j�  j/  j  Kj~  K�hhChAh`ubK�j�  )��}�(j�  KHj�  j�  j�  j1  j  Kj~  K�hhChAh�ubK�j�  )��}�(j�  KHj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  Kj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  KNj�  j�  j�  jE  j  K'j~  K�hhChAh�ubK�j�  )��}�(j�  KNj�  j�  j�  jG  j  K'j~  K�hhChAh�ubK�j�  )��}�(j�  KNj�  j�  j�  j  )��}�(h^j�  h>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  K'j~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  KOj�  j�  j�  j3  j  K(j~  K�hhChAh`ubK�j�  )��}�(j�  KOj�  j�  j�  j7  j  K(j~  K�hhChAhiubK�j�  )��}�(j�  KOj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  K
hj�~  hAj�~  ubj  K(j~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  KOj�  j�  j�  j5  j  K)j~  K�hhChAh`ubK�j�  )��}�(j�  KOj�  j�  j�  j9  j  K)j~  K�hhChAhiubK�j�  )��}�(j�  KOj�  j�  j�  jC  j  K)j~  K�hh�hAh�ubK�j�  )��}�(j�  KOj�  j�  j�  j;  j  K*j~  K�hhChAh`ubK�j�  )��}�(j�  KOj�  j�  j�  j?  j  K*j~  K�hhChAhiubK�j�  )��}�(j�  KOj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  K*j~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  KNj�  j�  j�  j=  j  K*j~  K�hhChAh�ubK�j�  )��}�(j�  KNj�  j�  j�  jA  j  K*j~  K�hhChAh�ubK�j�  )��}�(j�  KNj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  K*j~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  KFj�  j�  j�  j[  j  K6j~  K�hhChAhqubK�j�  )��}�(j�  KFj�  j�  j�  jU  j  K6j~  K�hhChAh�ubK�j�  )��}�(j�  KFj�  j�  j�  jW  j  K6j~  K�hh�hAh�ubK�j�  )��}�(j�  KFj�  j�  j�  j[  j  K6j~  K�hhChAhqubK�j�  )��}�(j�  KFj�  j�  j�  jY  j  K6j~  K�hhChAhfubK�j�  )��}�(j�  KFj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  K6j~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  KFj�  j�  j�  j[  j  K6j~  K�hhChAhqubK�j�  )��}�(j�  KFj�  j�  j�  j]  j  K6j~  K�hhChAhfubK�j�  )��}�(j�  KFj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  K	hj�~  hAj�~  ubj  K6j~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  K/j�  j�  j�  jl  j  KKj~  K�hhChAh`ubK�j�  )��}�(j�  K/j�  j�  j�  jc  j  KKj~  K�hhChAhiubK�j�  )��}�(j�  K/j�  j�  j�  jg  j  KKj~  K�hji  hAjk  ubK�j�  )��}�(j�  K/j�  j�  j�  jl  j  KKj~  K�hhChAh`ubK�j�  )��}�(j�  K/j�  j�  j�  jt  j  KKj~  K�hhChAhfubK�j�  )��}�(j�  K/j�  j�  j�  jx  j  KKj~  K�hh�hAh�ubK�j�  )��}�(j�  K/j�  j�  j�  jn  j  KLj~  K�hhChAh`ubK�j�  )��}�(j�  K/j�  j�  j�  jr  j  KLj~  K�hhChAhNubK�j�  )��}�(j�  K/j�  j�  j�  jp  j  KMj~  K�hhChAh`ubK�j�  )��}�(j�  K/j�  j�  j�  jv  j  KMj~  K�hhChAhNubK�j�  )��}�(j�  KCj�  j�  j�  j|  j  KRj~  K�hhChAhqubK�j�  )��}�(j�  KCj�  j�  j�  jz  j  KRj~  K�hhChAh�ubK�j�  )��}�(j�  KCj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  KRj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  KCj�  j�  j�  j|  j  KRj~  K�hhChAhqubK�j�  )��}�(j�  KCj�  j�  j�  hb)��}�(h=KhKh>heh^ji�  hDhEhF�hG�h<�h_KhhChAhfubj  KRj~  K�hhChAhfubK�j�  )��}�(j�  KCj�  j�  j�  j  )��}�(h^jm�  h>h<hDj�~  hG�h<�j�~  K
hj�~  hAj�~  ubj  KRj~  K�hj�~  hAj�~  ubK�j�  )��}�(j�  KFj�  j�  j�  h)��}�(h=KhKh>h]h^NhDhEhF�hG�h<�h_KhhChAh�ubj  KRj~  K�hhChAh�ubK�j�  )��}�(j�  KFj�  j�  j�  j~  j  KRj~  K�hhChAh�ubK�j�  )��}�(j�  KFj�  j�  j�  j  )��}�(h^Nh>h<hDj�~  hG�h<�j�~  Khj�~  hAj�~  ubj  KRj~  K�hj�~  hAj�~  ubK�j�  K�j�  )��}�(j�  KFj�  j�  j�  hZ)��}�(h=KhKh>h]h^j{�  hDhEhF�hG�h<�h_K
hhChAh`ubj  KRj~  K�hhChAh`ubK�j�  )��}�(j�  KFj�  j�  j�  hs)��}�(h^j�  h<�h-Kh=Kh>hvh@�hKhAhrhB�hKhhChDhEhF�hG�hKhHKubj  KRj~  K�hhChAhrubu�args�]�(KKe�	equipList�]�(j�|  j  j�|  hzhshOh�hjh�h�hhbhZj�|  hnh�j  e�	tilesSeen�]��inSeed�J�x �cLevel�Kubj�  h	j  KRj~  KFhAhubj�~  Nj�~  K hD]�(KKYK�e�rightScroll�N�healthCurve�G?�333333j�~  K�Class��Player_Classes��
Spellsword���heh�)��}�(h=KhKh>hehDhEhF�hG�h<�h_KhhChAh�ubh]hZ)��}�(h=KhKh>h]hDhEhF�hG�h<�h_K
hhChAh`ubub�width�K#�turn�M{	j�  j�  �xConst�K�yConst�KF�MessageHandler�j�  �height�K�console��tdl��Console���)��K_K/]�(K K K K ��K K K ����KGK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KLK�K�K���K K K ����KEK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KRK�K�K���K K K ����KPK�K�K���K K K ����KAK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KWK�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KxK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KaK�K�K���K K K ����KoK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KFK�K�K���K K K ����K K K K ��K K K ����KvK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KnK�K�K���K K K ����KwK�K�K���K K K ����KmK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KoK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KoK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KoK�K�K���K K K ����KbK�K�K���K K K ����KoK�K�K���K K K ����KbK�K�K���K K K ����KoK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KwK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KgK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KgK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KgK�K�K���K K K ����KiK�K�K���K K K ����KgK�K�K���K K K ����KiK�K�K���K K K ����KgK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K1K�K�K���K K K ����K K K K ��K K K ����KhK�K�K���K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K:K�K�K���K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KPK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K1K�K�K���K K K ����K5K�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KpK�K�K���K K K ����KAK�K�K���K K K ����KAK�K�K���K K K ����KaK�K�K���K K K ����KAK�K�K���K K K ����KAK�K�K���K K K ����KAK�K�K���K K K ����KAK�K�K���K K K ����KAK�K�K���K K K ����KGK�K�K���K K K ����KpK�K�K���K K K ����KGK�K�K���K K K ����KaK�K�K���K K K ����KGK�K�K���K K K ����KaK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K4K�K�K���K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K9K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KiK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KtK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KiK�K�K���K K K ����KrK�K�K���K K K ����KcK�K�K���K K K ����KrK�K�K���K K K ����KtK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KAK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K9K�K�K���K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KtK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KuK�K�K���K K K ����KcK�K�K���K K K ����KuK�K�K���K K K ����KqK�K�K���K K K ����KuK�K�K���K K K ����KtK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K9K�K�K���K K K ����K K K K ��K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KkK�K�K���K K K ����KhK�K�K���K K K ����KhK�K�K���K K K ����KaK�K�K���K K K ����KhK�K�K���K K K ����KhK�K�K���K K K ����KhK�K�K���K K K ����KhK�K�K���K K K ����KhK�K�K���K K K ����KnK�K�K���K K K ����KkK�K�K���K K K ����KnK�K�K���K K K ����KuK�K�K���K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KcK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KtK�K�K���K K K ����KeK�K�K���K K K ����KtK�K�K���K K K ����KiK�K�K���K K K ����KtK�K�K���K K K ����KcK�K�K���K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KSK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K �����       K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KdK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KkK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K�K�K���K K K ����KdK�K�K���K K K ����K K�K�K���K K K ����KrK�K�K���K K K ����K K�K�K���K K K ����KkK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KpK�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����KmK�K�K���K K K ����KeK�K�K���K K K ����KiK�K�K���K K K ����KwK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KcK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KuK�K�K���K K K ����KaK�K�K���K K K ����KaK�K�K���K K K ����KdK�K�K���K K K ����KiK�K�K���K K K ����KwK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KiK�K�K���K K K ����KuK�K�K���K K K ����KtK�K�K���K K K ����KdK�K�K���K K K ����KiK�K�K���K K K ����KdK�K�K���K K K ����KsK�K�K���K K K ����KaK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KkK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KpK�K�K���K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����KaK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KcK�K�K���K K K ����KpK�K�K���K K K ����KtK�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����KGK�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KkK�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����K5K�K�K���K K K ����KsK�K�K���K K K ����KGK�K�K���K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KIK�K�K���K K K ����KaK�K�K���K K K ����KaK�K�K���K K K ����KoK�K�K���K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KeK�K�K���K K K ����KBK�K�K���K K K ����KcK�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����KfK�K�K���K K K ����KkK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KrK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KbK�K�K���K K K ����KfK�K�K���K K K ����KkK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KdK�K�K���K K K ����KoK�K�K���K K K ����KkK�K�K���K K K ����KcK�K�K���K K K ����KdK�K�K���K K K ����KbK�K�K���K K K ����KrK�K�K���K K K ����KiK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KTK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KoK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KlK�K�K���K K K ����KrK�K�K���K K K ����KiK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����KwK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����KlK�K�K���K K K ����KaK�K�K���K K K ����KlK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KiK�K�K���K K K ����KaK�K�K���K K K ����KlK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KuK�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����KiK�K�K���K K K ����KGK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KwK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KnK�K�K���K K K ����KiK�K�K���K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����KnK�K�K���K K K ����KdK�K�K���K K K ����KeK�K�K���K K K ����KBK�K�K���K K K ����KLK�K�K���K K K ����KLK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KHK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KdK�K�K���K K K ����KeK�K�K���K K K ����KCK�K�K���K K K ����KBK�K�K���K K K ����KGK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����KsK�K�K���K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����K!K�K�K���K K K ����KdK�K�K���K K K ����KuK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KGK�K�K���K K K ����KGK�K�K���K K K ����KAK�K�K���K K K ����K!K�K�K���K K K ����KdK�K�K���K K K ����KlK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KCK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KcK�K�K���K K K ����KaK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KlK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KoK�K�K���K K K ����KwK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KbK�K�K���K K K ����KkK�K�K���K K K ����KtK�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����KmK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KcK�K�K���K K K ����K K K K ��K K K ����KbK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KuK�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����KlK�K�K���K K K ����KhK�K�K���K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KwK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KgK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KCK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KrK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KfK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KfK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����KdK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����KfK�K�K���K K K ����KfK�K�K���K K K ����KfK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KsK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K4K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K1K�K�K���K K K ����K4K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����e(K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K$K�K�K��K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K@KKYK���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K?K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K=KQKOK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K4K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KSK�K�K���K K K ����KLK�K�K���K K K ����KRK�K�K���K K K ����KDK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KFK�K�K���K K K ����KLK�K�K���K K K ����KRK�K�K���K K K ����KDK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KLK�K�K���K K K ����KLK�K�K���K K K ����KRK�K�K���K K K ����KDK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KhK�K�K���K K K ����KeK�K�K���K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KeK�K�K���K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KeK�K�K���K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KvK�K�K���K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KvK�K�K���K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KvK�K�K���K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KcK�K�K���K K K ����KeK�K�K���K K K ����KgK�K�K���K K K ����KlK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KgK�K�K���K K K ����KlK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KhK�K�K���K K K ����KeK�K�K���K K K ����KgK�K�K���K K K ����KlK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KkK�K�K���K K K ����KlK�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����KbK�K�K���K K K ����KlK�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KlK�K�K���K K K ����KeK�K�K���K K K ����KsK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KmK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K1K�K�K���K K K ����K1K�K�K���K K K ����KiK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K1K�K�K���K K K ����K5K�K�K���K K K ����KaK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K1K�K�K���K K K ����K5K�K�K���K K K ����KmK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KfK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KcK�K�K���K K K ����KuK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KfK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����KBK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KcK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KmK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KcK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KpK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KcK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����KcK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ���[0      K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KcK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e��bub.