��      �Player�h ��)��}�(�	sightDist�K�accuracy�K �	rightHand��Items.Weapons��Staff���)��}�(�armorPen�K�level�K�range�K�color�]�(K�K�K�e�type��2H��
equippable���addPower���magPower�K�
usesArrows���char��?��weight�K�	throwable���power�K�name��Staff��
consumable��ubhK�visible���canMove���arrows�K �invertColor��h�@��skillLevels�}�(�6�K �2�K �3�K �7�K �1�K �5�K �4�K u�gold�K hK�armorVal�K hK �rightScroll�N�skillPoints�KhK�
baseHealth�K��skills�}�(h&�	Abilities��Flash_Freeze���h'h4�Shocking_Grasp���h(h4�Fireball���h)h4�Arcane_Reservoir���h*h4�Blink���h+h4�Wall_of_Force���h,h4�Lightning_Bolt���u�
healthTemp�K �	rightRing�N�playerControlled���expNext�Kd�healthCurve�G?�      �	healthMax�K�h�Kyle��dodge�K �Class��Player_Classes��Mage����items�]�(�Items.Consumables��	GreenHerb���)��}�(�healNum�Kh�h�h�+�hhh�
Green Herb�h�
consumable�ubhS)��}�(hVKh�h�hhWhhhhXhhYube�
initiative�K�effects�]�h]�(KKYK�e�exp�K �
leftScroll�N�recalcTimer�K �leftRing�N�
hitEffects�]��helmet��Items.Armors��	Cloth_Hat���)��}�(h�h�hKhhhKh.Kh�hhh�	Cloth Hat�h�helmet�ub�health�K��
countering���	recalcMax�K �pObject��Object�hr��)��}�(�row�K"�ID�Khh#�pLevel��LevelTypes.LevelTypes��Wild���)��}�(�	decorList�]�(�LevelTypes.Decorations��Table���h��Firepit���h��Weapon_Rack���e�	thePlayer�h�master_Changed_Tiles�]�(]�(K!K@e]�(K K?e]�(KK>e]�(KK=e]�(KK<e]�(KK;e]�(KK:e]�(KK9e]�(K!KBe]�(K KCe]�(K!K@e]�(K K?e]�(KK>e]�(KK=e]�(KK<e]�(KK;e]�(KK:e]�(KK9e]�(K!KBe]�(K KCe]�(K!K@e]�(K K?e]�(KK>e]�(KK=e]�(KK<e]�(KK;e]�(KK:e]�(KK9e]�(K!KBe]�(K KCe]�(K!K@e]�(K K?e]�(K K>e]�(KK=e]�(KK<e]�(KK;e]�(KK:e]�(KK9e]�(K!KBe]�(K!KCe]�(K!K@e]�(K!K?e]�(K!KBe]�(K!KCe]�(K!K@e]�(K!K?e]�(K!KBe]�(K!KCe]�(K!K@e]�(K!K?e]�(K"KBe]�(K!KCe]�(K"K@e]�(K!K?e]�(K"KBe]�(K!KCe]�(K"K@e]�(K!K?e]�(K"KBe]�(K!KCe]�(K"K@e]�(K!K?e]�(K"KBe]�(K"KCe]�(K"K@e]�(K"K?e]�(K!K>e]�(K!K=e]�(K!K<e]�(K!K;e]�(K!K:e]�(K"KBe]�(K"KCe]�(K"K@e]�(K"K?e]�(K"K>e]�(K"K=e]�(K"K<e]�(K!K;e]�(K!K:e]�(K"KBe]�(K"KCe]�(K"K@e]�(K"K?e]�(K"K>e]�(K"K=e]�(K"K<e]�(K"K;e]�(K"K:e]�(K"KBe]�(K"KCe]�(K"K@e]�(K"K?e]�(K"K>e]�(K"K=e]�(K"K<e]�(K#K;e]�(K#K:e]�(K"KBe]�(K"KCe]�(K"K@e]�(K"K?e]�(K#K>e]�(K#K=e]�(K#K<e]�(K#K;e]�(K#K:e]�(K"KBe]�(K"KCe]�(K"K@e]�(K#K?e]�(K#K>e]�(K#K=e]�(K#K<e]�(K$K;e]�(K$K:e]�(K"KBe]�(K"KCe]�(K"K@e]�(K#K?e]�(K#K>e]�(K#K=e]�(K$K<e]�(K$K;e]�(K$K:e]�(K"KBe]�(K#KCe]�(K"K@e]�(K#K?e]�(K#K>e]�(K$K=e]�(K$K<e]�(K%K;e]�(K%K:e]�(K%K9e]�(K"KBe]�(K#KCe]�(K#K@e]�(K#K?e]�(K$K>e]�(K$K=e]�(K%K<e]�(K%K;e]�(K&K:e]�(K"KBe]�(K#KCe]�(K#K@e]�(K#K?e]�(K$K>e]�(K$K=e]�(K%K<e]�(K&K;e]�(K&K:e]�(K#KBe]�(K#KCe]�(K#K@e]�(K#K?e]�(K$K>e]�(K%K=e]�(K%K<e]�(K&K;e]�(K'K:e]�(K'K9e]�(K#KBe]�(K#KCe]�(K#K@e]�(K$K?e]�(K$K>e]�(K%K=e]�(K&K<e]�(K'K;e]�(K'K:e]�(K(K9e]�(K#KBe]�(K#KCe]�(K#K@e]�(K$K?e]�(K%K>e]�(K%K=e]�(K&K<e]�(K'K;e]�(K(K:e]�(K)K9e]�(K#KBe]�(K$KCe]�(K#K@e]�(K$K?e]�(K%K>e]�(K&K=e]�(K#KBe]�(K$KCe]�(K#K@e]�(K$K?e]�(K%K>e]�(K&K=e]�(K#KBe]�(K$KCe]�(K!K@e]�(K K?e]�(KK>e]�(KK=e]�(KK<e]�(KK;e]�(KK:e]�(KK9e]�(K#K@e]�(K$K?e]�(K%K>e]�(K&K=e]�(K!K@e]�(K K?e]�(KK>e]�(KK=e]�(KK<e]�(KK;e]�(KK;e]�(K#K@e]�(K$K?e]�(K%K>e]�(K&K=e]�(K!K@e]�(K K?e]�(KK>e]�(KK>e]�(KK=e]�(KK<e]�(KK;e]�(K#K@e]�(K$K?e]�(K%K?e]�(K&K>e]�(K!K@e]�(K K?e]�(KK?e]�(KK>e]�(KK=e]�(KK<e]�(KK<e]�(KK;e]�(K#K@e]�(K$K@e]�(K!K@e]�(K K@e]�(K#K@e]�(K$K@e]�(K!K@e]�(K K@e]�(K#K@e]�(K$K@e]�(K!K@e]�(K K@e]�(K#KAe]�(K$K@e]�(K!KAe]�(K#KAe]�(K$K@e]�(K!KAe]�(K#KAe]�(K$K@e]�(K!KAe]�(K#KAe]�(K$KAe]�(K%K@e]�(K&K@e]�(K'K@e]�(K(K@e]�(K)K?e]�(K*K?e]�(K!KAe]�(K#KAe]�(K$KAe]�(K%KAe]�(K&K@e]�(K'K@e]�(K(K@e]�(K)K@e]�(K*K@e]�(K!KAe]�(K#KAe]�(K$KAe]�(K%KAe]�(K&KAe]�(K'KAe]�(K(KAe]�(K)K@e]�(K*K@e]�(K!KAe]�(K#KAe]�(K$KAe]�(K%KAe]�(K&KAe]�(K'KAe]�(K(KAe]�(K)KAe]�(K*KAe]�(K!KAe]�(K#KAe]�(K$KAe]�(K%KAe]�(K&KAe]�(K'KAe]�(K(KAe]�(K)KBe]�(K*KBe]�(K!KAe]�(K#KAe]�(K$KAe]�(K%KAe]�(K&KBe]�(K'KBe]�(K(KBe]�(K)KBe]�(K*KBe]�(K!KAe]�(K#KAe]�(K$KAe]�(K%KBe]�(K&KBe]�(K'KBe]�(K(KBe]�(K)KCe]�(K!KAe]�(K#KAe]�(K$KBe]�(K%KBe]�(K&KBe]�(K'KCe]�(K!KAe]�(K#KAe]�(K$KBe]�(K%KBe]�(K&KCe]�(K!KBe]�(K KBe]�(KKCe]�(K#KAe]�(K$KBe]�(K%KBe]�(K&KCe]�(K!KBe]�(K KBe]�(KKCe]�(K#KBe]�(K$KBe]�(K%KCe]�(K!KBe]�(K KBe]�(KKCe]�(K#KBe]�(K$KBe]�(K%KCe]�(K!KBe]�(K KCe]�(K#KBe]�(K$KBe]�(K%KCe]�(K!KBe]�(K KCe]�(K#KBe]�(K$KCe]�(K!KBe]�(K KCe]�(K#KBe]�(K$KCe]�(K!KBe]�(K KCe]�(K#KBe]�(K$KCee�
stairsDown�]�(KAK"e�Tiles�}�(K }�(K �Tile�j�  ��)��}�(hvK �Objects�]�hxh|�col�K ubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubK	j   )��}�(hvK j  ]�hxh|j  K	ubK
j   )��}�(hvK j  ]�hxh|j  K
ubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubK j   )��}�(hvK j  ]�hxh|j  K ubK!j   )��}�(hvK j  ]�hxh|j  K!ubK"j   )��}�(hvK j  ]�hxh|j  K"ubK#j   )��}�(hvK j  ]�hxh|j  K#ubK$j   )��}�(hvK j  ]�hxh|j  K$ubK%j   )��}�(hvK j  ]�hxh|j  K%ubK&j   )��}�(hvK j  ]�hxh|j  K&ubK'j   )��}�(hvK j  ]�hxh|j  K'ubK(j   )��}�(hvK j  ]�hxh|j  K(ubK)j   )��}�(hvK j  ]�hxh|j  K)ubK*j   )��}�(hvK j  ]�hxh|j  K*ubK+j   )��}�(hvK j  ]�hxh|j  K+ubK,j   )��}�(hvK j  ]�hxh|j  K,ubK-j   )��}�(hvK j  ]�hxh|j  K-ubK.j   )��}�(hvK j  ]�hxh|j  K.ubK/j   )��}�(hvK j  ]�hxh|j  K/ubK0j   )��}�(hvK j  ]�hxh|j  K0ubK1j   )��}�(hvK j  ]�hxh|j  K1ubK2j   )��}�(hvK j  ]�hxh|j  K2ubK3j   )��}�(hvK j  ]�hxh|j  K3ubK4j   )��}�(hvK j  ]�hxh|j  K4ubK5j   )��}�(hvK j  ]�hxh|j  K5ubK6j   )��}�(hvK j  ]�hxh|j  K6ubK7j   )��}�(hvK j  ]�hxh|j  K7ubK8j   )��}�(hvK j  ]�hxh|j  K8ubK9j   )��}�(hvK j  ]�hxh|j  K9ubK:j   )��}�(hvK j  ]�hxh|j  K:ubK;j   )��}�(hvK j  ]�hxh|j  K;ubK<j   )��}�(hvK j  ]�hxh|j  K<ubK=j   )��}�(hvK j  ]�hxh|j  K=ubK>j   )��}�(hvK j  ]�hxh|j  K>ubK?j   )��}�(hvK j  ]�hxh|j  K?ubK@j   )��}�(hvK j  ]�hxh|j  K@ubKAj   )��}�(hvK j  ]�hxh|j  KAubKBj   )��}�(hvK j  ]�hxh|j  KBubKCj   )��}�(hvK j  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�K ahxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�Kahxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�Kahxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK	}�(K j   )��}�(hvK	j  ]�hxh|j  K ubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubK	j   )��}�(hvK	j  ]�hxh|j  K	ubK
j   )��}�(hvK	j  ]�hxh|j  K
ubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubKj   )��}�(hvK	j  ]�hxh|j  KubK j   )��}�(hvK	j  ]�hxh|j  K ubK!j   )��}�(hvK	j  ]�hxh|j  K!ubK"j   )��}�(hvK	j  ]�hxh|j  K"ubK#j   )��}�(hvK	j  ]�hxh|j  K#ubK$j   )��}�(hvK	j  ]�hxh|j  K$ubK%j   )��}�(hvK	j  ]�hxh|j  K%ubK&j   )��}�(hvK	j  ]�hxh|j  K&ubK'j   )��}�(hvK	j  ]�hxh|j  K'ubK(j   )��}�(hvK	j  ]�hxh|j  K(ubK)j   )��}�(hvK	j  ]�hxh|j  K)ubK*j   )��}�(hvK	j  ]�hxh|j  K*ubK+j   )��}�(hvK	j  ]�hxh|j  K+ubK,j   )��}�(hvK	j  ]�hxh|j  K,ubK-j   )��}�(hvK	j  ]�hxh|j  K-ubK.j   )��}�(hvK	j  ]�hxh|j  K.ubK/j   )��}�(hvK	j  ]�hxh|j  K/ubK0j   )��}�(hvK	j  ]�hxh|j  K0ubK1j   )��}�(hvK	j  ]�hxh|j  K1ubK2j   )��}�(hvK	j  ]�hxh|j  K2ubK3j   )��}�(hvK	j  ]�hxh|j  K3ubK4j   )��}�(hvK	j  ]�hxh|j  K4ubK5j   )��}�(hvK	j  ]�hxh|j  K5ubK6j   )��}�(hvK	j  ]�hxh|j  K6ubK7j   )��}�(hvK	j  ]�hxh|j  K7ubK8j   )��}�(hvK	j  ]�hxh|j  K8ubK9j   )��}�(hvK	j  ]�hxh|j  K9ubK:j   )��}�(hvK	j  ]�hxh|j  K:ubK;j   )��}�(hvK	j  ]�hxh|j  K;ubK<j   )��}�(hvK	j  ]�hxh|j  K<ubK=j   )��}�(hvK	j  ]�hxh|j  K=ubK>j   )��}�(hvK	j  ]�hxh|j  K>ubK?j   )��}�(hvK	j  ]�hxh|j  K?ubK@j   )��}�(hvK	j  ]�hxh|j  K@ubKAj   )��}�(hvK	j  ]�hxh|j  KAubKBj   )��}�(hvK	j  ]�hxh|j  KBubKCj   )��}�(hvK	j  ]�hxh|j  KCubuK
}�(K j   )��}�(hvK
j  ]�hxh|j  K ubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubK	j   )��}�(hvK
j  ]�hxh|j  K	ubK
j   )��}�(hvK
j  ]�hxh|j  K
ubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubKj   )��}�(hvK
j  ]�hxh|j  KubK j   )��}�(hvK
j  ]�hxh|j  K ubK!j   )��}�(hvK
j  ]�hxh|j  K!ubK"j   )��}�(hvK
j  ]�hxh|j  K"ubK#j   )��}�(hvK
j  ]�hxh|j  K#ubK$j   )��}�(hvK
j  ]�hxh|j  K$ubK%j   )��}�(hvK
j  ]�hxh|j  K%ubK&j   )��}�(hvK
j  ]�hxh|j  K&ubK'j   )��}�(hvK
j  ]�hxh|j  K'ubK(j   )��}�(hvK
j  ]�hxh|j  K(ubK)j   )��}�(hvK
j  ]�hxh|j  K)ubK*j   )��}�(hvK
j  ]�hxh|j  K*ubK+j   )��}�(hvK
j  ]�hxh|j  K+ubK,j   )��}�(hvK
j  ]�hxh|j  K,ubK-j   )��}�(hvK
j  ]�hxh|j  K-ubK.j   )��}�(hvK
j  ]�hxh|j  K.ubK/j   )��}�(hvK
j  ]�hxh|j  K/ubK0j   )��}�(hvK
j  ]�hxh|j  K0ubK1j   )��}�(hvK
j  ]�hxh|j  K1ubK2j   )��}�(hvK
j  ]�hxh|j  K2ubK3j   )��}�(hvK
j  ]�hxh|j  K3ubK4j   )��}�(hvK
j  ]�hxh|j  K4ubK5j   )��}�(hvK
j  ]�hxh|j  K5ubK6j   )��}�(hvK
j  ]�hxh|j  K6ubK7j   )��}�(hvK
j  ]�hxh|j  K7ubK8j   )��}�(hvK
j  ]�hxh|j  K8ubK9j   )��}�(hvK
j  ]�hxh|j  K9ubK:j   )��}�(hvK
j  ]�hxh|j  K:ubK;j   )��}�(hvK
j  ]�hxh|j  K;ubK<j   )��}�(hvK
j  ]�hxh|j  K<ubK=j   )��}�(hvK
j  ]�hxh|j  K=ubK>j   )��}�(hvK
j  ]�hxh|j  K>ubK?j   )��}�(hvK
j  ]�hxh|j  K?ubK@j   )��}�(hvK
j  ]�hxh|j  K@ubKAj   )��}�(hvK
j  ]�hxh|j  KAubKBj   )��}�(hvK
j  ]�hxh|j  KBubKCj   )��}�(hvK
j  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�Kahxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�Kahxh|j  K5ubK6j   )��}�(hvKj  ]�Kahxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  �       KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�Kahxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�Kahxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�Kahxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�hxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�K	ahxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�hxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK}�(K j   )��}�(hvKj  ]�hxh|j  K ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK	j   )��}�(hvKj  ]�hxh|j  K	ubK
j   )��}�(hvKj  ]�hxh|j  K
ubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubKj   )��}�(hvKj  ]�hxh|j  KubK j   )��}�(hvKj  ]�hxh|j  K ubK!j   )��}�(hvKj  ]�hxh|j  K!ubK"j   )��}�(hvKj  ]�hxh|j  K"ubK#j   )��}�(hvKj  ]�K
ahxh|j  K#ubK$j   )��}�(hvKj  ]�hxh|j  K$ubK%j   )��}�(hvKj  ]�hxh|j  K%ubK&j   )��}�(hvKj  ]�hxh|j  K&ubK'j   )��}�(hvKj  ]�hxh|j  K'ubK(j   )��}�(hvKj  ]�hxh|j  K(ubK)j   )��}�(hvKj  ]�hxh|j  K)ubK*j   )��}�(hvKj  ]�hxh|j  K*ubK+j   )��}�(hvKj  ]�hxh|j  K+ubK,j   )��}�(hvKj  ]�hxh|j  K,ubK-j   )��}�(hvKj  ]�hxh|j  K-ubK.j   )��}�(hvKj  ]�Kahxh|j  K.ubK/j   )��}�(hvKj  ]�hxh|j  K/ubK0j   )��}�(hvKj  ]�hxh|j  K0ubK1j   )��}�(hvKj  ]�hxh|j  K1ubK2j   )��}�(hvKj  ]�hxh|j  K2ubK3j   )��}�(hvKj  ]�hxh|j  K3ubK4j   )��}�(hvKj  ]�hxh|j  K4ubK5j   )��}�(hvKj  ]�hxh|j  K5ubK6j   )��}�(hvKj  ]�hxh|j  K6ubK7j   )��}�(hvKj  ]�hxh|j  K7ubK8j   )��}�(hvKj  ]�hxh|j  K8ubK9j   )��}�(hvKj  ]�hxh|j  K9ubK:j   )��}�(hvKj  ]�hxh|j  K:ubK;j   )��}�(hvKj  ]�hxh|j  K;ubK<j   )��}�(hvKj  ]�hxh|j  K<ubK=j   )��}�(hvKj  ]�hxh|j  K=ubK>j   )��}�(hvKj  ]�hxh|j  K>ubK?j   )��}�(hvKj  ]�hxh|j  K?ubK@j   )��}�(hvKj  ]�hxh|j  K@ubKAj   )��}�(hvKj  ]�hxh|j  KAubKBj   )��}�(hvKj  ]�hxh|j  KBubKCj   )��}�(hvKj  ]�hxh|j  KCubuK }�(K j   )��}�(hvK j  ]�hxh|j  K ubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubK	j   )��}�(hvK j  ]�hxh|j  K	ubK
j   )��}�(hvK j  ]�hxh|j  K
ubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubKj   )��}�(hvK j  ]�hxh|j  KubK j   )��}�(hvK j  ]�hxh|j  K ubK!j   )��}�(hvK j  ]�hxh|j  K!ubK"j   )��}�(hvK j  ]�hxh|j  K"ubK#j   )��}�(hvK j  ]�hxh|j  K#ubK$j   )��}�(hvK j  ]�hxh|j  K$ubK%j   )��}�(hvK j  ]�hxh|j  K%ubK&j   )��}�(hvK j  ]�hxh|j  K&ubK'j   )��}�(hvK j  ]�hxh|j  K'ubK(j   )��}�(hvK j  ]�hxh|j  K(ubK)j   )��}�(hvK j  ]�hxh|j  K)ubK*j   )��}�(hvK j  ]�hxh|j  K*ubK+j   )��}�(hvK j  ]�hxh|j  K+ubK,j   )��}�(hvK j  ]�hxh|j  K,ubK-j   )��}�(hvK j  ]�hxh|j  K-ubK.j   )��}�(hvK j  ]�hxh|j  K.ubK/j   )��}�(hvK j  ]�hxh|j  K/ubK0j   )��}�(hvK j  ]�hxh|j  K0ubK1j   )��}�(hvK j  ]�hxh|j  K1ubK2j   )��}�(hvK j  ]�hxh|j  K2ubK3j   )��}�(hvK j  ]�hxh|j  K3ubK4j   )��}�(hvK j  ]�hxh|j  K4ubK5j   )��}�(hvK j  ]�hxh|j  K5ubK6j   )��}�(hvK j  ]�hxh|j  K6ubK7j   )��}�(hvK j  ]�hxh|j  K7ubK8j   )��}�(hvK j  ]�hxh|j  K8ubK9j   )��}�(hvK j  ]�hxh|j  K9ubK:j   )��}�(hvK j  ]�hxh|j  K:ubK;j   )��}�(hvK j  ]�hxh|j  K;ubK<j   )��}�(hvK j  ]�hxh|j  K<ubK=j   )��}�(hvK j  ]�hxh|j  K=ubK>j   )��}�(hvK j  ]�hxh|j  K>ubK?j   )��}�(hvK j  ]�hxh|j  K?ubK@j   )��}�(hvK j  ]�hxh|j  K@ubKAj   )��}�(hvK j  ]�hxh|j  KAubKBj   )��}�(hvK j  ]�hxh|j  KBubKCj   )��}�(hvK j  ]�hxh|j  KCubuK!}�(K j   )��}�(hvK!j  ]�hxh|j  K ubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubK	j   )��}�(hvK!j  ]�hxh|j  K	ubK
j   )��}�(hvK!j  ]�hxh|j  K
ubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubKj   )��}�(hvK!j  ]�hxh|j  KubK j   )��}�(hvK!j  ]�hxh|j  K ubK!j   )��}�(hvK!j  ]�hxh|j  K!ubK"j   )��}�(hvK!j  ]�hxh|j  K"ubK#j   )��}�(hvK!j  ]�hxh|j  K#ubK$j   )��}�(hvK!j  ]�hxh|j  K$ubK%j   )��}�(hvK!j  ]�hxh|j  K%ubK&j   )��}�(hvK!j  ]�hxh|j  K&ubK'j   )��}�(hvK!j  ]�hxh|j  K'ubK(j   )��}�(hvK!j  ]�hxh|j  K(ubK)j   )��}�(hvK!j  ]�hxh|j  K)ubK*j   )��}�(hvK!j  ]�hxh|j  K*ubK+j   )��}�(hvK!j  ]�hxh|j  K+ubK,j   )��}�(hvK!j  ]�hxh|j  K,ubK-j   )��}�(hvK!j  ]�hxh|j  K-ubK.j   )��}�(hvK!j  ]�hxh|j  K.ubK/j   )��}�(hvK!j  ]�hxh|j  K/ubK0j   )��}�(hvK!j  ]�hxh|j  K0ubK1j   )��}�(hvK!j  ]�hxh|j  K1ubK2j   )��}�(hvK!j  ]�hxh|j  K2ubK3j   )��}�(hvK!j  ]�hxh|j  K3ubK4j   )��}�(hvK!j  ]�hxh|j  K4ubK5j   )��}�(hvK!j  ]�hxh|j  K5ubK6j   )��}�(hvK!j  ]�hxh|j  K6ubK7j   )��}�(hvK!j  ]�hxh|j  K7ubK8j   )��}�(hvK!j  ]�hxh|j  K8ubK9j   )��}�(hvK!j  ]�hxh|j  K9ubK:j   )��}�(hvK!j  ]�hxh|j  K:ubK;j   )��}�(hvK!j  ]�hxh|j  K;ubK<j   )��}�(hvK!j  ]�hxh|j  K<ubK=j   )��}�(hvK!j  ]�hxh|j  K=ubK>j   )��}�(hvK!j  ]�hxh|j  K>ubK?j   )��}�(hvK!j  ]�hxh|j  K?ubK@j   )��}�(hvK!j  ]�hxh|j  K@ubKAj   )��}�(hvK!j  ]�hxh|j  KAubKBj   )��}�(hvK!j  ]�hxh|j  KBubKCj   )��}�(hvK!j  ]�hxh|j  KCubuK"}�(K j   )��}�(hvK"j  ]�hxh|j  K ubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubK	j   )��}�(hvK"j  ]�hxh|j  K	ubK
j   )��}�(hvK"j  ]�hxh|j  K
ubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubKj   )��}�(hvK"j  ]�hxh|j  KubK j   )��}�(hvK"j  ]�hxh|j  K ubK!j   )��}�(hvK"j  ]�hxh|j  K!ubK"j   )��}�(hvK"j  ]�hxh|j  K"ubK#j   )��}�(hvK"j  ]�hxh|j  K#ubK$j   )��}�(hvK"j  ]�hxh|j  K$ubK%j   )��}�(hvK"j  ]�hxh|j  K%ubK&j   )��}�(hvK"j  ]�hxh|j  K&ubK'j   )��}�(hvK"j  ]�hxh|j  K'ubK(j   )��}�(hvK"j  ]�hxh|j  K(ubK)j   )��}�(hvK"j  ]�hxh|j  K)ubK*j   )��}�(hvK"j  ]�hxh|j  K*ubK+j   )��}�(hvK"j  ]�hxh|j  K+ubK,j   )��}�(hvK"j  ]�hxh|j  K,ubK-j   )��}�(hvK"j  ]�hxh|j  K-ubK.j   )��}�(hvK"j  ]�hxh|j  K.ubK/j   )��}�(hvK"j  ]�hxh|j  K/ubK0j   )��}�(hvK"j  ]�hxh|j  K0ubK1j   )��}�(hvK"j  ]�hxh|j  K1ubK2j   )��}�(hvK"j  ]�hxh|j  K2ubK3j   )��}�(hvK"j  ]�hxh|j  K3ubK4j   )��}�(hvK"j  ]�hxh|j  K4ubK5j   )��}�(hvK"j  ]�hxh|j  K5ubK6j   )��}�(hvK"j  ]�hxh|j  K6ubK7j   )��}�(hvK"j  ]�hxh|j  K7ubK8j   )��}�(hvK"j  ]�hxh|j  K8ubK9j   )��}�(hvK"j  ]�hxh|j  K9ubK:j   )��}�(hvK"j  ]�hxh|j  K:ubK;j   )��}�(hvK"j  ]�hxh|j  K;ubK<j   )��}�(hvK"j  ]�hxh|j  K<ubK=j   )��}�(hvK"j  ]�hxh|j  K=ubK>j   )��}�(hvK"j  ]�hxh|j  K>ubK?j   )��}�(hvK"j  ]�hxh|j  K?ubK@j   )��}�(hvK"j  ]�hxh|j  K@ubKAj   )��}�(hvK"j  ]�(KKehxh|j  KAubKBj   )��}�(hvK"j  ]�hxh|j  KBubKCj   )��}�(hvK"j  ]�hxh|j  KCubuK#}�(K j   )��}�(hvK#j  ]�hxh|j  K ubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubK	j   )��}�(hvK#j  ]�hxh|j  K	ubK
j   )��}�(hvK#j  ]�hxh|j  K
ubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubKj   )��}�(hvK#j  ]�hxh|j  KubK j   )��}�(hvK#j  ]�hxh|j  K ubK!j   )��}�(hvK#j  ]�hxh|j  K!ubK"j   )��}�(hvK#j  ]�hxh|j  K"ubK#j   )��}�(hvK#j  ]�hxh|j  K#ubK$j   )��}�(hvK#j  ]�hxh|j  K$ubK%j   )��}�(hvK#j  ]�hxh|j  K%ubK&j   )��}�(hvK#j  ]�hxh|j  K&ubK'j   )��}�(hvK#j  ]�hxh|j  K'ubK(j   )��}�(hvK#j  ]�hxh|j  K(ubK)j   )��}�(hvK#j  ]�hxh|j  K)ubK*j   )��}�(hvK#j  ]�hxh|j  K*ubK+j   )��}�(hvK#j  ]�hxh|j  K+ubK,j   )��}�(hvK#j  ]�hxh|j  K,ubK-j   )��}�(hvK#j  ]�hxh|j  K-ubK.j   )��}�(hvK#j  ]�hxh|j  K.ubK/j   )��}�(hvK#j  ]�hxh|j  K/ubK0j   )��}�(hvK#j  ]�hxh|j  K0ubK1j   )��}�(hvK#j  ]�hxh|j  K1ubK2j   )��}�(hvK#j  ]�hxh|j  K2ubK3j   )��}�(hvK#j  ]�hxh|j  K3ubK4j   )��}�(hvK#j  ]�hxh|j  K4ubK5j   )��}�(hvK#j  ]�hxh|j  K5ubK6j   )��}�(hvK#j  ]�hxh|j  K6ubK7j   )��}�(hvK#j  ]�hxh|j  K7ubK8j   )��}�(hvK#j  ]�hxh|j  K8ubK9j   )��}�(hvK#j  ]�hxh|j  K9ubK:j   )��}�(hvK#j  ]�hxh|j  K:ubK;j   )��}�(hvK#j  ]�hxh|j  K;ubK<j   )��}�(hvK#j  ]�hxh|j  K<ubK=j   )��}�(hvK#j  ]�hxh|j  K=ubK>j   )��}�(hvK#j  ]�hxh|j  K>ubK?j   )��}�(hvK#j  ]�hxh|j  K?ubK@j   )��}�(hvK#j  ]�hxh|j  K@ubKAj   )��}�(hvK#j  ]�hxh|j  KAubKBj   )��}�(hvK#j  ]�hxh|j  KBubKCj   )��}�(hvK#j  ]�hxh|j  KCubuK$}�(K j   )��}�(hvK$j  ]�hxh|j  K ubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubK	j   )��}�(hvK$j  ]�hxh|j  K	ubK
j   )��}�(hvK$j  ]�hxh|j  K
ubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubKj   )��}�(hvK$j  ]�hxh|j  KubK j   )��}�(hvK$j  ]�hxh|j  K ubK!j   )��}�(hvK$j  ]�hxh|j  K!ubK"j   )��}�(hvK$j  ]�hxh|j  K"ubK#j   )��}�(hvK$j  ]�hxh|j  K#ubK$j   )��}�(hvK$j  ]�hxh|j  K$ubK%j   )��}�(hvK$j  ]�hxh|j  K%ubK&j   )��}�(hvK$j  ]�hxh|j  K&ubK'j   )��}�(hvK$j  ]�hxh|j  K'ubK(j   )��}�(hvK$j  ]�hxh|j  K(ubK)j   )��}�(hvK$j  ]�hxh|j  K)ubK*j   )��}�(hvK$j  ]�hxh|j  K*ubK+j   )��}�(hvK$j  ]�hxh|j  K+ubK,j   )��}�(hvK$j  ]�hxh|j  K,ubK-j   )��}�(hvK$j  ]�hxh|j  K-ubK.j   )��}�(hvK$j  ]�hxh|j  K.ubK/j   )��}�(hvK$j  ]�hxh|j  K/ubK0j   )��}�(hvK$j  ]�hxh|j  K0ubK1j   )��}�(hvK$j  ]�hxh|j  K1ubK2j   )��}�(hvK$j  ]�hxh|j  K2ubK3j   )��}�(hvK$j  ]�hxh|j  K3ubK4j   )��}�(hvK$j  ]�hxh|j  K4ubK5j   )��}�(hvK$j  ]�hxh|j  K5ubK6j   )��}�(hvK$j  ]�hxh|j  K6ubK7j   )��}�(hvK$j  ]�hxh|j  K7ubK8j   )��}�(hvK$j  ]�hxh|j  K8ubK9j   )��}�(hvK$j  ]�hxh|j  K9ubK:j   )��}�(hvK$j  ]�hxh|j  K:ubK;j   )��}�(hvK$j  ]�hxh|j  K;ubK<j   )��}�(hvK$j  ]�hxh|j  K<ubK=j   )��}�(hvK$j  ]�hxh|j  K=ubK>j   )��}�(hvK$j  ]�hxh|j  K>ubK?j   )��}�(hvK$j  ]�hxh|j  K?ubK@j   )��}�(hvK$j  ]�hxh|j  K@ubKAj   )��}�(hvK$j  ]�hxh|j  KAubKBj   )��}�(hvK$j  ]�hxh|j  KBubKCj   )��}�(hvK$j  ]�hxh|j  KCubuK%}�(K j   )��}�(hvK%j  ]�hxh|j  K ubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubK	j   )��}�(hvK%j  ]�hxh|j  K	ubK
j   )��}�(hvK%j  ]�hxh|j  K
ubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubKj   )��}�(hvK%j  ]�hxh|j  KubK j   )��}�(hvK%j  ]�hxh|j  K ubK!j   )��}�(hvK%j  ]�hxh|j  K!ubK"j   )��}�(hvK%j  ]�hxh|j  K"ubK#j   )��}�(hvK%j  ]�hxh|j  K#ubK$j   )��}�(hvK%j  ]�hxh|j  K$ubK%j   )��}�(hvK%j  ]�hxh|j  K%ubK&j   )��}�(hvK%j  ]�hxh|j  K&ubK'j   )��}�(hvK%j  ]�hxh|j  K'ubK(j   )��}�(hvK%j  ]�hxh|j  K(ubK)j   )��}�(hvK%j  ]�hxh|j  K)ubK*j   )��}�(hvK%j  ]�hxh|j  K*ubK+j   )��}�(hvK%j  ]�hxh|j  K+ubK,j   )��}�(hvK%j  ]�hxh|j  K,ubK-j   )��}�(hvK%j  ]�hxh|j  K-ubK.j   )��}�(hvK%j  ]�hxh|j  K.ubK/j   )��}�(hvK%j  ]�hxh|j  K/ubK0j   )��}�(hvK%j  ]�hxh|j  K0ubK1j   )��}�(hvK%j  ]�hxh|j  K1ubK2j   )��}�(hvK%j  ]�hxh|j  K2ubK3j   )��}�(hvK%j  ]�hxh|j  K3ubK4j   )��}�(hvK%j  ]�hxh|j  K4ubK5j   )��}�(hvK%j  ]�hxh|j  K5ubK6j   )��}�(hvK%j  ]�hxh|j  K6ubK7j   )��}�(hvK%j  ]�hxh|j  K7ubK8j   )��}�(hvK%j  ]�hxh|j  K8ubK9j   )��}�(hvK%j  ]�hxh|j  K9ubK:j   )��}�(hvK%j  ]�hxh|j  K:ubK;j   )��}�(hvK%j  ]�hxh|j  K;ubK<j   )��}�(hvK%j  ]�hxh|j  K<ubK=j   )��}�(hvK%j  ]�hxh|j  K=ubK>j   )��}�(hvK%j  ]�hxh|j  K>ubK?j   )��}�(hvK%j  ]�hxh|j  K?ubK@j   )��}�(hvK%j  ]�hxh|j  K@ubKAj   )��}�(hvK%j  ]�hxh|j  KAubKBj   )��}�(hvK%j  ]�hxh|j  KBubKCj   )��}�(hvK%j  ]�hxh|j  KCubuK&}�(K j   )��}�(hvK&j  ]�hxh|j  K ubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubK	j   )��}�(hvK&j  ]�hxh|j  K	ubK
j   )��}�(hvK&j  ]�hxh|j  K
ubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubKj   )��}�(hvK&j  ]�hxh|j  KubK j   )��}�(hvK&j  ]�hxh|j  K ubK!j   )��}�(hvK&j  ]�hxh|j  K!ubK"j   )��}�(hvK&j  ]�hxh|j  K"ubK#j   )��}�(hvK&j  ]�hxh|j  K#ubK$j   )��}�(hvK&j  ]�hxh|j  K$ubK%j   )��}�(hvK&j  ]�hxh|j  K%ubK&j   )��}�(hvK&j  ]�hxh|j  K&ubK'j   )��}�(hvK&j  ]�hxh|j  K'ubK(j   )��}�(hvK&j  ]�hxh|j  K(ubK)j   )��}�(hvK&j  ]�hxh|j  K)ubK*j   )��}�(hvK&j  ]�hxh|j  K*ubK+j   )��}�(hvK&j  ]�hxh|j  K+ubK,j   )��}�(hvK&j  ]�hxh|j  K,ubK-j   )��}�(hvK&j  ]�hxh|j  K-ubK.j   )��}�(hvK&j  ]�hxh|j  K.ubK/j   )��}�(hvK&j  ]�hxh|j  K/ubK0j   )��}�(hvK&j  ]�hxh|j  K0ubK1j   )��}�(hvK&j  ]�hxh|j  K1ubK2j   )��}�(hvK&j  ]�hxh|j  K2ubK3j   )��}�(hvK&j  ]�hxh|j  K3ubK4j   )��}�(hvK&j  ]�hxh|j  K4ubK5j   )��}�(hvK&j  ]�hxh|j  K5ubK6j   )��}�(hvK&j  ]�hxh|j  K6ubK7j   )��}�(hvK&j  ]�hxh|j  K7ubK8j   )��}�(hvK&j  ]�hxh|j  K8ubK9j   )��}�(hvK&j  ]�hxh|j  K9ubK:j   )��}�(hvK&j  ]�hxh|j  K:ubK;j   )��}�(hvK&j  ]�hxh|j  K;ubK<j   )��}�(hvK&j  ]�hxh|j  K<ubK=j   )��}�(hvK&j  ]�hxh|j  K=ubK>j   )��}�(hvK&j  ]�hxh|j  K>ubK?j   )��}�(hvK&j  ]�hxh|j  K?ubK@j   )��}�(hvK&j  ]�hxh|j  K@ubKAj   )��}�(hvK&j  ]�hxh|j  KAubKBj   )��}�(hvK&j  ]�hxh|j  KBubKCj   )��}�(hvK&j  ]�hxh|j  KCubuK'}�(K j   )��}�(hvK'j  ]�hxh|j  K ubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubK	j   )��}�(hvK'j  ]�hxh|j  K	ubK
j   )��}�(hvK'j  ]�hxh|j  K
ubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubKj   )��}�(hvK'j  ]�hxh|j  KubK j   )��}�(hvK'j  ]�hxh|j  K ubK!j   )��}�(hvK'j  ]�hxh|j  K!ubK"j   )��}�(hvK'j  ]�hxh|j  K"ubK#j   )��}�(hvK'j  ]�hxh|j  K#ubK$j   )��}�(hvK'j  ]�hxh|j  K$ubK%j   )��}�(hvK'j  ]�hxh|j  K%ubK&j   )��}�(hvK'j  ]�hxh|j  K&ubK'j   )��}�(hvK'j  ]�hxh|j  K'ubK(j   )��}�(hvK'j  ]�hxh|j  K(ubK)j   )��}�(hvK'j  ]�hxh|j  K)ubK*j   )��}�(hvK'j  ]�hxh|j  K*ubK+j   )��}�(hvK'j  ]�hxh|j  K+ubK,j   )��}�(hvK'j  ]�hxh|j  K,ubK-j   )��}�(hvK'j  ]�hxh|j  K-ubK.j   )��}�(hvK'j  ]�hxh|j  K.ubK/j   )��}�(hvK'j  ]�hxh|j  K/ubK0j   )��}�(hvK'j  ]�hxh|j  K0ubK1j   )��}�(hvK'j  ]�hxh|j  K1ubK2j   )��}�(hvK'j  ]�hxh|j  K2ubK3j   )��}�(hvK'j  ]�hxh|j  K3ubK4j   )��}�(hvK'j  ]�hxh|j  K4ubK5j   )��}�(hvK'j  ]�hxh|j  K5ubK6j   )��}�(hvK'j  ]�hxh|j  K6ubK7j   )��}�(hvK'j  ]�hxh|j  K7ubK8j   )��}�(hvK'j  ]�hxh|j  K8ubK9j   )��}�(hvK'j  ]�hxh|j  K9ubK:j   )��}�(hvK'j  ]�hxh|j  K:ubK;j   )��}�(hvK'j  ]�hxh|j  K;ubK<j   )��}�(hvK'j  ]�hxh|j  K<ubK=j   )��}�(hvK'j  ]�hxh|j  K=ubK>j   )��}�(hvK'j  ]�hxh|j  K>ubK?j   )��}�(hvK'j  ]�hxh|j  K?ubK@j   )��}�(hvK'j  ]�hxh|j  K@ubKAj   )��}�(hvK'j  ]�hxh|j  KAubKBj   )��}�(hvK'j  ]�hxh|j  KBubKCj   )��}�(hvK'j  ]�hxh|j  KCubuK(}�(K j   )��}�(hvK(j  ]�hxh|j  K ubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubK	j   )��}�(hvK(j  ]�hxh|j  K	ubK
j   )��}�(hvK(j  ]�hxh|j  K
ubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubKj   )��}�(hvK(j  ]�hxh|j  KubK j   )��}�(hvK(j  ]�hxh|j  K ubK!j   )��}�(hvK(j  ]�hxh|j  K!ubK"j   )��}�(hvK(j  ]�hxh|j  K"ubK#j   )��}�(hvK(j  ]�hxh|j  K#ubK$j   )��}�(hvK(j  ]�hxh|j  K$ubK%j   )��}�(hvK(j  ]�hxh|j  K%ubK&j   )��}�(hvK(j  ]�hxh|j  K&ubK'j   )��}�(hvK(j  ]�hxh|j  K'ubK(j   )��}�(hvK(j  ]�hxh|j  K(ubK)j   )��}�(hvK(j  ]�hxh|j  K)ubK*j   )��}�(hvK(j  ]�hxh|j  K*ubK+j   )��}�(hvK(j  ]�hxh|j  K+ubK,j   )��}�(hvK(j  ]�hxh|j  K,ubK-j   )��}�(hvK(j  ]�hxh|j  K-ubK.j   )��}�(hvK(j  ]�hxh|j  K.ubK/j   )��}�(hvK(j  ]�hxh|j  K/ubK0j   )��}�(hvK(j  ]�hxh|j  K0ubK1j   )��}�(hvK(j  ]�hxh|j  K1ubK2j   )��}�(hvK(j  ]�hxh|j  K2ubK3j   )��}�(hvK(j  ]�hxh|j  K3ubK4j   )��}�(hvK(j  ]�hxh|j  K4ubK5j   )��}�(hvK(j  ]�hxh|j  K5ubK6j   )��}�(hvK(j  ]�hxh|j  K6ubK7j   )��}�(hvK(j  ]�hxh|j  K7ubK8j   )��}�(hvK(j  ]�hxh|j  K8ubK9j   )��}�(hvK(j  ]�hxh|j  K9ubK:j   )��}�(hvK(j  ]�hxh|j  K:ubK;j   )��}�(hvK(j  ]�hxh|j  K;ubK<j   )��}�(hvK(j  ]�hxh|j  K<ubK=j   )��}�(hvK(j  ]�hxh|j  K=ubK>j   )��}�(hvK(j  ]�hxh|j  K>ubK?j   )��}�(hvK(j  ]�hxh|j  K?ubK@j   )��}�(hvK(j  ]�hxh|j  K@ubKAj   )��}�(hvK(j  ]�hxh|j  KAubKBj   )��}�(hvK(j  ]�hxh|j  KBubKCj   )��}�(hvK(j  ]�hxh|j  KCubuK)}�(K j   )��}�(hvK)j  ]�hxh|j  K ubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubK	j   )��}�(hvK)j  ]�hxh|j  K	ubK
j   )��}�(hvK)j  ]�hxh|j  K
ubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubKj   )��}�(hvK)j  ]�hxh|j  KubK j   )��}�(hvK)j  ]�hxh|j  K ubK!j   )��}�(hvK)j  ]�hxh|j  K!ubK"j   )��}�(hvK)j  ]�hxh|j  K"ubK#j   )��}�(hvK)j  ]�hxh|j  K#ubK$j   )��}�(hvK)j  ]�hxh|j  K$ubK%j   )��}�(hvK)j  ]�hxh|j  K%ubK&j   )��}�(hvK)j  ]�hxh|j  K&ubK'j   )��}�(hvK)j  ]�hxh|j  K'ubK(j   )��}�(hvK)j  ]�hxh|j  K(ubK)j   )��}�(hvK)j  ]�hxh|j  K)ubK*j   )��}�(hvK)j  ]�hxh|j  K*ubK+j   )��}�(hvK)j  ]�hxh|j  K+ubK,j   )��}�(hvK)j  ]�hxh|j  K,ubK-j   )��}�(hvK)j  ]�hxh|j  K-ubK.j   )��}�(hvK)j  ]�hxh|j  K.ubK/j   )��}�(hvK)j  ]�hxh|j  K/ubK0j   )��}�(hvK)j  ]�hxh|j  K0ubK1j   )��}�(hvK)j  ]�hxh|j  K1ubK2j   )��}�(hvK)j  ]�hxh|j  K2ubK3j   )��}�(hvK)j  ]�hxh|j  K3ubK4j   )��}�(hvK)j  ]�hxh|j  K4ubK5j   )��}�(hvK)j  ]�hxh|j  K5ubK6j   )��}�(hvK)j  ]�hxh|j  K6ubK7j   )��}�(hvK)j  ]�hxh|j  K7ubK8j   )��}�(hvK)j  ]�hxh|j  K8ubK9j   )��}�(hvK)j  ]�hxh|j  K9ubK:j   )��}�(hvK)j  ]�hxh|j  K:ubK;j   )��}�(hvK)j  ]�hxh|j  K;ubK<j   )��}�(hvK)j  ]�hxh|j  K<ubK=j   )��}�(hvK)j  ]�hxh|j  K=ubK>j   )��}�(hvK)j  ]�hxh|j  K>ubK?j   )��}�(hvK)j  ]�hxh|j  K?ubK@j   )��}�(hvK)j  ]�hxh|j  K@ubKAj   )��}�(hvK)j  ]�hxh|j  KAubKBj   )��}�(hvK)j  ]�hxh|j  KBubKCj   )��}�(hvK)j  ]�hxh|j  KCubuK*}�(K j   )��}�(hvK*j  ]�hxh|j  K ubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubK	j   )��}�(hvK*j  ]�hxh|j  K	ubK
j   )��}�(hvK*j  ]�hxh|j  K
ubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubKj   )��}�(hvK*j  ]�hxh|j  KubK j   )��}�(hvK*j  ]�hxh|j  K ubK!j   )��}�(hvK*j  ]�hxh|j  K!ubK"j   )��}�(hvK*j  ]�hxh|j  K"ubK#j   )��}�(hvK*j  ]�hxh|j  K#ubK$j   )��}�(hvK*j  ]�hxh|j  K$ubK%j   )��}�(hvK*j  ]�hxh|j  K%ubK&j   )��}�(hvK*j  ]�hxh|j  K&ubK'j   )��}�(hvK*j  ]�hxh|j  K'ubK(j   )��}�(hvK*j  ]�hxh|j  K(ubK)j   )��}�(hvK*j  ]�hxh|j  K)ubK*j   )��}�(hvK*j  ]�hxh|j  K*ubK+j   )��}�(hvK*j  ]�hxh|j  K+ubK,j   )��}�(hvK*j  ]�hxh|j  K,ubK-j   )��}�(hvK*j  ]�hxh|j  K-ubK.j   )��}�(hvK*j  ]�hxh|j  K.ubK/j   )��}�(hvK*j  ]�hxh|j  K/ubK0j   )��}�(hvK*j  ]�hxh|j  K0ubK1j   )��}�(hvK*j  ]�hxh|j  K1ubK2j   )��}�(hvK*j  ]�hxh|j  K2ubK3j   )��}�(hvK*j  ]�hxh|j  K3ubK4j   )��}�(hvK*j  ]�hxh|j  K4ubK5j   )��}�(hvK*j  ]�hxh|j  K5ubK6j   )��}�(hvK*j  ]�hxh|j  K6ubK7j   )��}�(hvK*j  ]�hxh|j  K7ubK8j   )��}�(hvK*j  ]�hxh|j  K8ubK9j   )��}�(hvK*j  ]�hxh|j  K9ubK:j   )��}�(hvK*j  ]�hxh|j  K:ubK;j   )��}�(hvK*j  ]�hxh|j  K;ubK<j   )��}�(hvK*j  ]�hxh|j  K<ubK=j   )��}�(hvK*j  ]�hxh|j  K=ubK>j   )��}�(hvK*j  ]�hxh|j  K>ubK?j   )��}�(hvK*j  ]�hxh|j  K?ubK@j   )��}�(hvK*j  ]�hxh|j  K@ubKAj   )��}�(hvK*j  ]�hxh|j  KAubKBj   )��}�(hvK*j  ]�hxh|j  KBubKCj   )��}�(hvK*j  ]�hxh|j  KCubuK+}�(K j   )��}�(hvK+j  ]�hxh|j  K ubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubK	j   )��}�(hvK+j  ]�hxh|j  K	ubK
j   )��}�(hvK+j  ]�hxh|j  K
ubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubKj   )��}�(hvK+j  ]�hxh|j  KubK j   )��}�(hvK+j  ]�hxh|j  K ubK!j   )��}�(hvK+j  ]�hxh|j  K!ubK"j   )��}�(hvK+j  ]�hxh|j  K"ubK#j   )��}�(hvK+j  ]�hxh|j  K#ubK$j   )��}�(hvK+j  ]�hxh|j  K$ubK%j   )��}�(hvK+j  ]�hxh|j  K%ubK&j   )��}�(hvK+j  ]�hxh|j  K&ubK'j   )��}�(hvK+j  ]�hxh|j  K'ubK(j   )��}�(hvK+j  ]�hxh|j  K(ubK)j   )��}�(hvK+j  ]�hxh|j  K)ubK*j   )��}�(hvK+j  ]�hxh|j  K*ubK+j   )��}�(hvK+j  ]�hxh|j  K+ubK,j   )��}�(hvK+j  ]�hxh|j  K,ubK-j   )��}�(hvK+j  ]�hxh|j  K-ubK.j   )��}�(hvK+j  ]�hxh|j  K.ubK/j   )��}�(hvK+j  ]�hxh|j  K/ubK0j   )��}�(hvK+j  ]�hxh|j  K0ubK1j   )��}�(hvK+j  ]�hxh|j  K1ubK2j   )��}�(hvK+j  ]�hxh|j  K2ubK3j   )��}�(hvK+j  ]�hxh|j  K3ubK4j   )��}�(hvK+j  ]�hxh|j  K4ubK5j   )��}�(hvK+j  ]�hxh|j  K5ubK6j   )��}�(hvK+j  ]�hxh|j  K6ubK7j   )��}�(hvK+j  ]�hxh|j  K7ubK8j   )��}�(hvK+j  ]�hxh|j  K8ubK9j   )��}�(hvK+j  ]�hxh|j  K9ubK:j   )��}�(hvK+j  ]�hxh|j  K:ubK;j   )��}�(hvK+j  ]�hxh|j  K;ubK<j   )��}�(hvK+j  ]�hxh|j  K<ubK=j   )��}�(hvK+j  ]�hxh|j  K=ubK>j   )��}�(hvK+j  ]�hxh|j  K>ubK?j   )��}�(hvK+j  ]�hxh|j  K?ubK@j   )��}�(hvK+j  ]�hxh|j  K@ubKAj   )��}�(hvK+j  ]�hxh|j  KAubKBj   )��}�(hvK+j  ]�hxh|j  KBubKCj   )��}�(hvK+j  ]�hxh|j  KCubuK,}�(K j   )��}�(hvK,j  ]�hxh|j  K ubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubK	j   )��}�(hvK,j  ]�hxh|j  K	ubK
j   )��}�(hvK,j  ]�hxh|j  K
ubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubKj   )��}�(hvK,j  ]�hxh|j  KubK j   )��}�(hvK,j  ]�hxh|j  K ubK!j   )��}�(hvK,j  ]�hxh|j  K!ubK"j   )��}�(hvK,j  ]�hxh|j  K"ubK#j   )��}�(hvK,j  ]�hxh|j  K#ubK$j   )��}�(hvK,j  ]�hxh|j  K$ubK%j   )��}�(hvK,j  ]�hxh|j  K%ubK&j   )��}�(hvK,j  ]�hxh|j  K&ubK'j   )��}�(hvK,j  ]�hxh|j  K'ubK(j   )��}�(hvK,j  ]�hxh|j  K(ubK)j   )��}�(hvK,j  ]�hxh|j  K)ubK*j   )��}�(hvK,j  ]�hxh|j  K*ubK+j   )��}�(hvK,j  ]�hxh|j  K+ubK,j   )��}�(hvK,j  ]�hxh|j  K,ubK-j   )��}�(hvK,j  ]�hxh|j  K-ubK.j   )��}�(hvK,j  ]�hxh|j  K.ubK/j   )��}�(hvK,j  ]�hxh|j  K/ubK0j   )��}�(hvK,j  ]�hxh|j  K0ubK1j   )��}�(hvK,j  ]�hxh|j  K1ubK2j   )��}�(hvK,j  ]�hxh|j  K2ubK3j   )��}�(hvK,j  ]�hxh|j  K3ubK4j   )��}�(hvK,j  ]�hxh|j  K4ubK5j   )��}�(hvK,j  ]�hxh|j  K5ubK6j   )��}�(hvK,j  ]�hxh|j  K6ubK7j   )��}�(hvK,j  ]�hxh|j  K7ubK8j   )��}�(hvK,j  ]�hxh|j  K8ubK9j   )��}�(hvK,j  ]�hxh|j  K9ubK:j   )��}�(hvK,j  ]�hxh|j  K:ubK;j   )��}�(hvK,j  ]�hxh|j  K;ubK<j   )��}�(hvK,j  ]�hxh|j  K<ubK=j   )��}�(hvK,j  ]�hxh|j  K=ubK>j   )��}�(hvK,j  ]�hxh|j  K>ubK?j   )��}�(hvK,j  ]�hxh|j  K?ubK@j   )��}�(hvK,j  ]�hxh|j  K@ubKAj   )��}�(hvK,j  ]�hxh|j  KAubKBj   )��}�(hvK,j  ]�hxh|j  KBubKCj   )��}�(hvK,j  ]�hxh|j  KCubuK-}�(K j   )��}�(hvK-j  ]�hxh|j  K ubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubK	j   )��}�(hvK-j  ]�hxh|j  K	ubK
j   )��}�(hvK-j  ]�hxh|j  K
ubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubKj   )��}�(hvK-j  ]�hxh|j  KubK j   )��}�(hvK-j  ]�hxh|j  K ubK!j   )��}�(hvK-j  ]�hxh|j  K!ubK"j   )��}�(hvK-j  ]�hxh|j  K"ubK#j   )��}�(hvK-j  ]�hxh|j  K#ubK$j   )��}�(hvK-j  ]�hxh|j  K$ubK%j   )��}�(hvK-j  ]�hxh|j  K%ubK&j   )��}�(hvK-j  ]�hxh|j  K&ubK'j   )��}�(hvK-j  ]�hxh|j  K'ubK(j   )��}�(hvK-j  ]�hxh|j  K(ubK)j   )��}�(hvK-j  ]�hxh|j  K)ubK*j   )��}�(hvK-j  ]�hxh|j  K*ubK+j   )��}�(hvK-j  ]�hxh|j  K+ubK,j   )��}�(hvK-j  ]�hxh|j  K,ubK-j   )��}�(hvK-j  ]�hxh|j  K-ubK.j   )��}�(hvK-j  ]�hxh|j  K.ubK/j   )��}�(hvK-j  ]�hxh|j  K/ubK0j   )��}�(hvK-j  ]�hxh|j  K0ubK1j   )��}�(hvK-j  ]�hxh|j  K1ubK2j   )��}�(hvK-j  ]�hxh|j  K2ubK3j   )��}�(hvK-j  ]�hxh|j  K3ubK4j   )��}�(hvK-j  ]�hxh|j  K4ubK5j   )��}�(hvK-j  ]�hxh|j  K5ubK6j   )��}�(hvK-j  ]�hxh|j  K6ubK7j   )��}�(hvK-j  ]�hxh|j  K7ubK8j   )��}�(hvK-j  ]�hxh|j  K8ubK9j   )��}�(hvK-j  ]�hxh|j  K9ubK:j   )��}�(hvK-j  ]�hxh|j  K:ubK;j   )��}�(hvK-j  ]�hxh|j  K;ubK<j   )��}�(hvK-j  ]�hxh|j  K<ubK=j   )��}�(hvK-j  ]�hxh|j  K=ubK>j   )��}�(hvK-j  ]�hxh|j  K>ubK?j   )��}�(hvK-j  ]�hxh|j  K?ubK@j   )��}�(hvK-j  ]�hxh|j  K@ubKAj   )��}�(hvK-j  ]�hxh|j  KAubKBj   )��}�(hvK-j  ]�hxh|j  KBubKCj   )��}�(hvK-j  ]�hxh|j  KCubuK.}�(K j   )��}�(hvK.j  ]�hxh|j  K ubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubK	j   )��}�(hvK.j  ]�hxh|j  K	ubK
j   )��}�(hvK.j  ]�hxh|j  K
ubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubKj   )��}�(hvK.j  ]�hxh|j  KubK j   )��}�(hvK.j  ]�hxh|j  K ubK!j   )��}�(hvK.j  ]�hxh|j  K!ubK"j   )��}�(hvK.j  ]�hxh|j  K"ubK#j   )��}�(hvK.j  ]�hxh|j  K#ubK$j   )��}�(hvK.j  ]�hxh|j  K$ubK%j   )��}�(hvK.j  ]�hxh|j  K%ubK&j   )��}�(hvK.j  ]�hxh|j  K&ubK'j   )��}�(hvK.j  ]�hxh|j  K'ubK(j   )��}�(hvK.j  ]�hxh|j  K(ubK)j   )��}�(hvK.j  ]�hxh|j  K)ubK*j   )��}�(hvK.j  ]�hxh|j  K*ubK+j   )��}�(hvK.j  ]�hxh|j  K+ubK,j   )��}�(hvK.j  ]�hxh|j  K,ubK-j   )��}�(hvK.j  ]�hxh|j  K-ubK.j   )��}�(hvK.j  ]�hxh|j  K.ubK/j   )��}�(hvK.j  ]�hxh|j  K/ubK0j   )��}�(hvK.j  ]�hxh|j  K0ubK1j   )��}�(hvK.j  ]�hxh|j  K1ubK2j   )��}�(hvK.j  ]�hxh|j  K2ubK3j   )��}�(hvK.j  ]�hxh|j  K3ubK4j   )��}�(hvK.j  ]�hxh|j  K4ubK5j   )��}�(hvK.j  ]�hxh|j  K5ubK6j   )��}�(hvK.j  ]�hxh|j  K6ubK7j   )��}�(hvK.j  ]�hxh|j  K7ubK8j   )��}�(hvK.j  ]�hxh|j  K8ubK9j   )��}�(hvK.j  ]�hxh|j  K9ubK:j   )��}�(hvK.j  ]�hxh|j  K:ubK;j   )��}�(hvK.j  ]�hxh|j  K;ubK<j   )��}�(hvK.j  ]�hxh|j  K<ubK=j   )��}�(hvK.j  ]�hxh|j  K=ubK>j   )��}�(hvK.j  ]�hxh|j  K>ubK?j   )��}�(hvK.j  ]�hxh|j  K?ubK@j   )��}�(hvK.j  ]�hxh|j  K@ubKAj   )��}�(hvK.j  ]�hxh|j  KAubKBj   )��}�(hvK.j  ]�hxh|j  KBubKCj   )��}�(hvK.j  ]�hxh|j  KCubuK/}�(K j   )��}�(hvK/j  ]�hxh|j  K ubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubK	j   )��}�(hvK/j  ]�hxh|j  K	ubK
j   )��}�(hvK/j  ]�hxh|j  K
ubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubKj   )��}�(hvK/j  ]�hxh|j  KubK j   )��}�(hvK/j  ]�hxh|j  K ubK!j   )��}�(hvK/j  ]�hxh|j  K!ubK"j   )��}�(hvK/j  ]�hxh|j  K"ubK#j   )��}�(hvK/j  ]�hxh|j  K#ubK$j   )��}�(hvK/j  ]�hxh|j  K$ubK%j   )��}�(hvK/j  ]�hxh|j  K%ubK&j   )��}�(hvK/j  ]�hxh|j  K&ubK'j   )��}�(hvK/j  ]�hxh|j  K'ubK(j   )��}�(hvK/j  ]�hxh|j  K(ubK)j   )��}�(hvK/j  ]�hxh|j  K)ubK*j   )��}�(hvK/j  ]�hxh|j  K*ubK+j   )��}�(hvK/j  ]�hxh|j  K+ubK,j   )��}�(hvK/j  ]�hxh|j  K,ubK-j   )��}�(hvK/j  ]�hxh|j  K-ubK.j   )��}�(hvK/j  ]�hxh|j  K.ubK/j   )��}�(hvK/j  ]�hxh|j  K/ubK0j   )��}�(hvK/j  ]�hxh|j  K0ubK1j   )��}�(hvK/j  ]�hxh|j  K1ubK2j   )��}�(hvK/j  ]�hxh|j  K2ubK3j   )��}�(hvK/j  ]�hxh|j  K3ubK4j   )��}�(hvK/j  ]�hxh|j  K4ubK5j   )��}�(hvK/j  ]�hxh|j  K5ubK6j   )��}�(hvK/j  ]�hxh|j  K6ubK7j   )��}�(hvK/j  ]�hxh|j  K7ubK8j   )��}�(hvK/j  ]�hxh|j  K8ubK9j   )��}�(hvK/j  ]�hxh|j  K9ubK:j   )��}�(hvK/j  ]�hxh|j  K:ubK;j   )��}�(hvK/j  ]�hxh|j  K;ubK<j   )��}�(hvK/j  ]�hxh|j  K<ubK=j   )��}�(hvK/j  ]�hxh|j  K=ubK>j   )��}�(hvK/j  ]�hxh|j  K>ubK?j   )��}�(hvK/j  ]�hxh|j  K?ubK@j   )��}�(hvK/j  ]�hxh|j  K@ubKAj   )��}�(hvK/j  ]�hxh|j  KAubKBj   )��}�(hvK/j  ]�hxh|j  KBubKCj   )��}�(hvK/j  ]�hxh|j  KCubuK0}�(K j   )��}�(hvK0j  ]�hxh|j  K ubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubK	j   )��}�(hvK0j  ]�hxh|j  K	ubK
j   )��}�(hvK0j  ]�hxh|j  K
ubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubKj   )��}�(hvK0j  ]�hxh|j  KubK j   )��}�(hvK0j  ]�hxh|j  K ubK!j   )��}�(hvK0j  ]�hxh|j  K!ubK"j   )��}�(hvK0j  ]�hxh|j  K"ubK#j   )��}�(hvK0j  ]�hxh|j  K#ubK$j   )��}�(hvK0j  ]�hxh|j  K$ubK%j   )��}�(hvK0j  ]�hxh|j  K%ubK&j   )��}�(hvK0j  ]�hxh|j  K&ubK'j   )��}�(hvK0j  ]�hxh|j  K'ubK(j   )��}�(hvK0j  ]�hxh|j  K(ubK)j   )��}�(hvK0j  ]�hxh|j  K)ubK*j   )��}�(hvK0j  ]�hxh|j  K*ubK+j   )��}�(hvK0j  ]�hxh|j  K+ubK,j   )��}�(hvK0j  ]�hxh|j  K,ubK-j   )��}�(hvK0j  ]�hxh|j  K-ubK.j   )��}�(hvK0j  ]�hxh|j  K.ubK/j   )��}�(hvK0j  ]�hxh|j  K/ubK0j   )��}�(hvK0j  ]�hxh|j  K0ubK1j   )��}�(hvK0j  ]�hxh|j  K1ubK2j   )��}�(hvK0j  ]�hxh|j  K2ubK3j   )��}�(hvK0j  ]�hxh|j  K3ubK4j   )��}�(hvK0j  ]�hxh|j  K4ubK5j   )��}�(hvK0j  ]�hxh|j  K5ubK6j   )��}�(hvK0j  ]�hxh|j  K6ubK7j   )��}�(hvK0j  ]�hxh|j  K7ubK8j   )��}�(hvK0j  ]�hxh|j  K8ubK9j   )��}�(hvK0j  ]�hxh|j  K9ubK:j   )��}�(hvK0j  ]�hxh|j  K:ubK;j   )��}�(hvK0j  ]�hxh|j  K;ubK<j   )��}�(hvK0j  ]�hxh|j  K<ubK=j   )��}�(hvK0j  ]�hxh|j  K=ubK>j   )��}�(hvK0j  ]�hxh|j  K>ubK?j   )��}�(hvK0j  ]�hxh|j  K?ubK@j   )��}�(hvK0j  ]�hxh|j  K@ubKAj   )��}�(hvK0j  ]�hxh|j  KAubKBj   )��}�(hvK0j  ]�hxh|j  KBubKCj   )��}�(hvK0j  ]�hxh|j  KCubuK1}�(K j   )��}�(hvK1j  ]�hxh|j  K ubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubK	j   )��}�(hvK1j  ]�hxh|j  K	ubK
j   )��}�(hvK1j  ]�hxh|j  K
ubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubKj   )��}�(hvK1j  ]�hxh|j  KubK j   )��}�(hvK1j  ]�hxh|j  K ubK!j   )��}�(hvK1j  ]�hxh|j  K!ubK"j   )��}�(hvK1j  ]�hxh|j  K"ubK#j   )��}�(hvK1j  ]�hxh|j  K#ubK$j   )��}�(hvK1j  ]�hxh|j  K$ubK%j   )��}�(hvK1j  ]�hxh|j  K%ubK&j   )��}�(hvK1j  ]�hxh|j  K&ubK'j   )��}�(hvK1j  ]�hxh|j  K'ubK(j   )��}�(hvK1j  ]�hxh|j  K(ubK)j   )��}�(hvK1j  ]�hxh|j  K)ubK*j   )��}�(hvK1j  ]�hxh|j  K*ubK+j   )��}�(hvK1j  ]�hxh|j  K+ubK,j   )��}�(hvK1j  ]�hxh|j  K,ubK-j   )��}�(hvK1j  ]�hxh|j  K-ubK.j   )��}�(hvK1j  ]�hxh|j  K.ubK/j   )��}�(hvK1j  ]�hxh|j  K/ubK0j   )��}�(hvK1j  ]�hxh|j  K0ubK1j   )��}�(hvK1j  ]�hxh|j  K1ubK2j   )��}�(hvK1j  ]�hxh|j  K2ubK3j   )��}�(hvK1j  ]�hxh|j  K3ubK4j   )��}�(hvK1j  ]�hxh|j  K4ubK5j   )��}�(hvK1j  ]�hxh|j  K5ubK6j   )��}�(hvK1j  ]�hxh|j  K6ubK7j   )��}�(hvK1j  ]�hxh|j  K7ubK8j   )��}�(hvK1j  ]�hxh|j  K8ubK9j   )��}�(hvK1j  ]�hxh|j  K9ubK:j   )��}�(hvK1j  ]�hxh|j  K:ubK;j   )��}�(hvK1j  ]�hxh|j  K;ubK<j   )��}�(hvK1j  ]�hxh|j  K<ubK=j   )��}�(hvK1j  ]�hxh|j  K=ubK>j   )��}�(hvK1j  ]�hxh|j  K>ubK?j   )��}�(hvK1j  ]�hxh|j  K?ubK@j   )��}�(hvK1j  ]�hxh|j  K@ubKAj   )��}�(hvK1j  ]�hxh|j  KAubKBj   )��}�(hvK1j  ]�hxh|j  KBubKCj   )��}�(hvK1j  ]�hxh|j  KCubuK2}�(K j   )��}�(hvK2j  ]�hxh|j  K ubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubK	j   )��}�(hvK2j  ]�hxh|j  K	ubK
j   )��}�(hvK2j  ]�hxh|j  K
ubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )���      }�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubKj   )��}�(hvK2j  ]�hxh|j  KubK j   )��}�(hvK2j  ]�hxh|j  K ubK!j   )��}�(hvK2j  ]�hxh|j  K!ubK"j   )��}�(hvK2j  ]�hxh|j  K"ubK#j   )��}�(hvK2j  ]�hxh|j  K#ubK$j   )��}�(hvK2j  ]�hxh|j  K$ubK%j   )��}�(hvK2j  ]�hxh|j  K%ubK&j   )��}�(hvK2j  ]�hxh|j  K&ubK'j   )��}�(hvK2j  ]�hxh|j  K'ubK(j   )��}�(hvK2j  ]�hxh|j  K(ubK)j   )��}�(hvK2j  ]�hxh|j  K)ubK*j   )��}�(hvK2j  ]�hxh|j  K*ubK+j   )��}�(hvK2j  ]�hxh|j  K+ubK,j   )��}�(hvK2j  ]�hxh|j  K,ubK-j   )��}�(hvK2j  ]�hxh|j  K-ubK.j   )��}�(hvK2j  ]�hxh|j  K.ubK/j   )��}�(hvK2j  ]�hxh|j  K/ubK0j   )��}�(hvK2j  ]�hxh|j  K0ubK1j   )��}�(hvK2j  ]�hxh|j  K1ubK2j   )��}�(hvK2j  ]�hxh|j  K2ubK3j   )��}�(hvK2j  ]�hxh|j  K3ubK4j   )��}�(hvK2j  ]�hxh|j  K4ubK5j   )��}�(hvK2j  ]�hxh|j  K5ubK6j   )��}�(hvK2j  ]�hxh|j  K6ubK7j   )��}�(hvK2j  ]�hxh|j  K7ubK8j   )��}�(hvK2j  ]�hxh|j  K8ubK9j   )��}�(hvK2j  ]�hxh|j  K9ubK:j   )��}�(hvK2j  ]�hxh|j  K:ubK;j   )��}�(hvK2j  ]�hxh|j  K;ubK<j   )��}�(hvK2j  ]�hxh|j  K<ubK=j   )��}�(hvK2j  ]�hxh|j  K=ubK>j   )��}�(hvK2j  ]�hxh|j  K>ubK?j   )��}�(hvK2j  ]�hxh|j  K?ubK@j   )��}�(hvK2j  ]�hxh|j  K@ubKAj   )��}�(hvK2j  ]�hxh|j  KAubKBj   )��}�(hvK2j  ]�hxh|j  KBubKCj   )��}�(hvK2j  ]�hxh|j  KCubuK3}�(K j   )��}�(hvK3j  ]�hxh|j  K ubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubK	j   )��}�(hvK3j  ]�hxh|j  K	ubK
j   )��}�(hvK3j  ]�hxh|j  K
ubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubKj   )��}�(hvK3j  ]�hxh|j  KubK j   )��}�(hvK3j  ]�hxh|j  K ubK!j   )��}�(hvK3j  ]�hxh|j  K!ubK"j   )��}�(hvK3j  ]�hxh|j  K"ubK#j   )��}�(hvK3j  ]�hxh|j  K#ubK$j   )��}�(hvK3j  ]�hxh|j  K$ubK%j   )��}�(hvK3j  ]�hxh|j  K%ubK&j   )��}�(hvK3j  ]�hxh|j  K&ubK'j   )��}�(hvK3j  ]�hxh|j  K'ubK(j   )��}�(hvK3j  ]�hxh|j  K(ubK)j   )��}�(hvK3j  ]�hxh|j  K)ubK*j   )��}�(hvK3j  ]�hxh|j  K*ubK+j   )��}�(hvK3j  ]�hxh|j  K+ubK,j   )��}�(hvK3j  ]�hxh|j  K,ubK-j   )��}�(hvK3j  ]�hxh|j  K-ubK.j   )��}�(hvK3j  ]�hxh|j  K.ubK/j   )��}�(hvK3j  ]�hxh|j  K/ubK0j   )��}�(hvK3j  ]�hxh|j  K0ubK1j   )��}�(hvK3j  ]�hxh|j  K1ubK2j   )��}�(hvK3j  ]�hxh|j  K2ubK3j   )��}�(hvK3j  ]�hxh|j  K3ubK4j   )��}�(hvK3j  ]�hxh|j  K4ubK5j   )��}�(hvK3j  ]�hxh|j  K5ubK6j   )��}�(hvK3j  ]�hxh|j  K6ubK7j   )��}�(hvK3j  ]�hxh|j  K7ubK8j   )��}�(hvK3j  ]�hxh|j  K8ubK9j   )��}�(hvK3j  ]�hxh|j  K9ubK:j   )��}�(hvK3j  ]�hxh|j  K:ubK;j   )��}�(hvK3j  ]�hxh|j  K;ubK<j   )��}�(hvK3j  ]�hxh|j  K<ubK=j   )��}�(hvK3j  ]�hxh|j  K=ubK>j   )��}�(hvK3j  ]�hxh|j  K>ubK?j   )��}�(hvK3j  ]�hxh|j  K?ubK@j   )��}�(hvK3j  ]�hxh|j  K@ubKAj   )��}�(hvK3j  ]�hxh|j  KAubKBj   )��}�(hvK3j  ]�hxh|j  KBubKCj   )��}�(hvK3j  ]�hxh|j  KCubuK4}�(K j   )��}�(hvK4j  ]�hxh|j  K ubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubK	j   )��}�(hvK4j  ]�hxh|j  K	ubK
j   )��}�(hvK4j  ]�hxh|j  K
ubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubKj   )��}�(hvK4j  ]�hxh|j  KubK j   )��}�(hvK4j  ]�hxh|j  K ubK!j   )��}�(hvK4j  ]�hxh|j  K!ubK"j   )��}�(hvK4j  ]�hxh|j  K"ubK#j   )��}�(hvK4j  ]�hxh|j  K#ubK$j   )��}�(hvK4j  ]�hxh|j  K$ubK%j   )��}�(hvK4j  ]�hxh|j  K%ubK&j   )��}�(hvK4j  ]�hxh|j  K&ubK'j   )��}�(hvK4j  ]�hxh|j  K'ubK(j   )��}�(hvK4j  ]�hxh|j  K(ubK)j   )��}�(hvK4j  ]�hxh|j  K)ubK*j   )��}�(hvK4j  ]�hxh|j  K*ubK+j   )��}�(hvK4j  ]�hxh|j  K+ubK,j   )��}�(hvK4j  ]�hxh|j  K,ubK-j   )��}�(hvK4j  ]�hxh|j  K-ubK.j   )��}�(hvK4j  ]�hxh|j  K.ubK/j   )��}�(hvK4j  ]�hxh|j  K/ubK0j   )��}�(hvK4j  ]�hxh|j  K0ubK1j   )��}�(hvK4j  ]�hxh|j  K1ubK2j   )��}�(hvK4j  ]�hxh|j  K2ubK3j   )��}�(hvK4j  ]�hxh|j  K3ubK4j   )��}�(hvK4j  ]�hxh|j  K4ubK5j   )��}�(hvK4j  ]�hxh|j  K5ubK6j   )��}�(hvK4j  ]�hxh|j  K6ubK7j   )��}�(hvK4j  ]�hxh|j  K7ubK8j   )��}�(hvK4j  ]�hxh|j  K8ubK9j   )��}�(hvK4j  ]�hxh|j  K9ubK:j   )��}�(hvK4j  ]�hxh|j  K:ubK;j   )��}�(hvK4j  ]�hxh|j  K;ubK<j   )��}�(hvK4j  ]�hxh|j  K<ubK=j   )��}�(hvK4j  ]�hxh|j  K=ubK>j   )��}�(hvK4j  ]�hxh|j  K>ubK?j   )��}�(hvK4j  ]�hxh|j  K?ubK@j   )��}�(hvK4j  ]�hxh|j  K@ubKAj   )��}�(hvK4j  ]�hxh|j  KAubKBj   )��}�(hvK4j  ]�hxh|j  KBubKCj   )��}�(hvK4j  ]�hxh|j  KCubuK5}�(K j   )��}�(hvK5j  ]�hxh|j  K ubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubK	j   )��}�(hvK5j  ]�hxh|j  K	ubK
j   )��}�(hvK5j  ]�hxh|j  K
ubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubKj   )��}�(hvK5j  ]�hxh|j  KubK j   )��}�(hvK5j  ]�hxh|j  K ubK!j   )��}�(hvK5j  ]�hxh|j  K!ubK"j   )��}�(hvK5j  ]�hxh|j  K"ubK#j   )��}�(hvK5j  ]�hxh|j  K#ubK$j   )��}�(hvK5j  ]�hxh|j  K$ubK%j   )��}�(hvK5j  ]�hxh|j  K%ubK&j   )��}�(hvK5j  ]�hxh|j  K&ubK'j   )��}�(hvK5j  ]�hxh|j  K'ubK(j   )��}�(hvK5j  ]�hxh|j  K(ubK)j   )��}�(hvK5j  ]�hxh|j  K)ubK*j   )��}�(hvK5j  ]�hxh|j  K*ubK+j   )��}�(hvK5j  ]�hxh|j  K+ubK,j   )��}�(hvK5j  ]�hxh|j  K,ubK-j   )��}�(hvK5j  ]�hxh|j  K-ubK.j   )��}�(hvK5j  ]�hxh|j  K.ubK/j   )��}�(hvK5j  ]�hxh|j  K/ubK0j   )��}�(hvK5j  ]�hxh|j  K0ubK1j   )��}�(hvK5j  ]�hxh|j  K1ubK2j   )��}�(hvK5j  ]�hxh|j  K2ubK3j   )��}�(hvK5j  ]�hxh|j  K3ubK4j   )��}�(hvK5j  ]�hxh|j  K4ubK5j   )��}�(hvK5j  ]�hxh|j  K5ubK6j   )��}�(hvK5j  ]�hxh|j  K6ubK7j   )��}�(hvK5j  ]�hxh|j  K7ubK8j   )��}�(hvK5j  ]�hxh|j  K8ubK9j   )��}�(hvK5j  ]�hxh|j  K9ubK:j   )��}�(hvK5j  ]�hxh|j  K:ubK;j   )��}�(hvK5j  ]�hxh|j  K;ubK<j   )��}�(hvK5j  ]�hxh|j  K<ubK=j   )��}�(hvK5j  ]�Kahxh|j  K=ubK>j   )��}�(hvK5j  ]�hxh|j  K>ubK?j   )��}�(hvK5j  ]�hxh|j  K?ubK@j   )��}�(hvK5j  ]�hxh|j  K@ubKAj   )��}�(hvK5j  ]�hxh|j  KAubKBj   )��}�(hvK5j  ]�hxh|j  KBubKCj   )��}�(hvK5j  ]�hxh|j  KCubuK6}�(K j   )��}�(hvK6j  ]�hxh|j  K ubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubK	j   )��}�(hvK6j  ]�hxh|j  K	ubK
j   )��}�(hvK6j  ]�hxh|j  K
ubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubKj   )��}�(hvK6j  ]�hxh|j  KubK j   )��}�(hvK6j  ]�hxh|j  K ubK!j   )��}�(hvK6j  ]�hxh|j  K!ubK"j   )��}�(hvK6j  ]�hxh|j  K"ubK#j   )��}�(hvK6j  ]�hxh|j  K#ubK$j   )��}�(hvK6j  ]�hxh|j  K$ubK%j   )��}�(hvK6j  ]�hxh|j  K%ubK&j   )��}�(hvK6j  ]�hxh|j  K&ubK'j   )��}�(hvK6j  ]�hxh|j  K'ubK(j   )��}�(hvK6j  ]�hxh|j  K(ubK)j   )��}�(hvK6j  ]�hxh|j  K)ubK*j   )��}�(hvK6j  ]�hxh|j  K*ubK+j   )��}�(hvK6j  ]�hxh|j  K+ubK,j   )��}�(hvK6j  ]�hxh|j  K,ubK-j   )��}�(hvK6j  ]�hxh|j  K-ubK.j   )��}�(hvK6j  ]�hxh|j  K.ubK/j   )��}�(hvK6j  ]�hxh|j  K/ubK0j   )��}�(hvK6j  ]�hxh|j  K0ubK1j   )��}�(hvK6j  ]�hxh|j  K1ubK2j   )��}�(hvK6j  ]�hxh|j  K2ubK3j   )��}�(hvK6j  ]�hxh|j  K3ubK4j   )��}�(hvK6j  ]�hxh|j  K4ubK5j   )��}�(hvK6j  ]�hxh|j  K5ubK6j   )��}�(hvK6j  ]�hxh|j  K6ubK7j   )��}�(hvK6j  ]�hxh|j  K7ubK8j   )��}�(hvK6j  ]�hxh|j  K8ubK9j   )��}�(hvK6j  ]�hxh|j  K9ubK:j   )��}�(hvK6j  ]�hxh|j  K:ubK;j   )��}�(hvK6j  ]�hxh|j  K;ubK<j   )��}�(hvK6j  ]�hxh|j  K<ubK=j   )��}�(hvK6j  ]�hxh|j  K=ubK>j   )��}�(hvK6j  ]�hxh|j  K>ubK?j   )��}�(hvK6j  ]�hxh|j  K?ubK@j   )��}�(hvK6j  ]�hxh|j  K@ubKAj   )��}�(hvK6j  ]�hxh|j  KAubKBj   )��}�(hvK6j  ]�hxh|j  KBubKCj   )��}�(hvK6j  ]�hxh|j  KCubuK7}�(K j   )��}�(hvK7j  ]�hxh|j  K ubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubK	j   )��}�(hvK7j  ]�hxh|j  K	ubK
j   )��}�(hvK7j  ]�hxh|j  K
ubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubKj   )��}�(hvK7j  ]�hxh|j  KubK j   )��}�(hvK7j  ]�hxh|j  K ubK!j   )��}�(hvK7j  ]�hxh|j  K!ubK"j   )��}�(hvK7j  ]�hxh|j  K"ubK#j   )��}�(hvK7j  ]�hxh|j  K#ubK$j   )��}�(hvK7j  ]�hxh|j  K$ubK%j   )��}�(hvK7j  ]�hxh|j  K%ubK&j   )��}�(hvK7j  ]�hxh|j  K&ubK'j   )��}�(hvK7j  ]�hxh|j  K'ubK(j   )��}�(hvK7j  ]�hxh|j  K(ubK)j   )��}�(hvK7j  ]�hxh|j  K)ubK*j   )��}�(hvK7j  ]�hxh|j  K*ubK+j   )��}�(hvK7j  ]�hxh|j  K+ubK,j   )��}�(hvK7j  ]�hxh|j  K,ubK-j   )��}�(hvK7j  ]�hxh|j  K-ubK.j   )��}�(hvK7j  ]�hxh|j  K.ubK/j   )��}�(hvK7j  ]�hxh|j  K/ubK0j   )��}�(hvK7j  ]�hxh|j  K0ubK1j   )��}�(hvK7j  ]�hxh|j  K1ubK2j   )��}�(hvK7j  ]�hxh|j  K2ubK3j   )��}�(hvK7j  ]�hxh|j  K3ubK4j   )��}�(hvK7j  ]�hxh|j  K4ubK5j   )��}�(hvK7j  ]�hxh|j  K5ubK6j   )��}�(hvK7j  ]�hxh|j  K6ubK7j   )��}�(hvK7j  ]�hxh|j  K7ubK8j   )��}�(hvK7j  ]�hxh|j  K8ubK9j   )��}�(hvK7j  ]�hxh|j  K9ubK:j   )��}�(hvK7j  ]�hxh|j  K:ubK;j   )��}�(hvK7j  ]�hxh|j  K;ubK<j   )��}�(hvK7j  ]�hxh|j  K<ubK=j   )��}�(hvK7j  ]�Kahxh|j  K=ubK>j   )��}�(hvK7j  ]�hxh|j  K>ubK?j   )��}�(hvK7j  ]�hxh|j  K?ubK@j   )��}�(hvK7j  ]�Kahxh|j  K@ubKAj   )��}�(hvK7j  ]�hxh|j  KAubKBj   )��}�(hvK7j  ]�hxh|j  KBubKCj   )��}�(hvK7j  ]�hxh|j  KCubuK8}�(K j   )��}�(hvK8j  ]�hxh|j  K ubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubK	j   )��}�(hvK8j  ]�hxh|j  K	ubK
j   )��}�(hvK8j  ]�hxh|j  K
ubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubKj   )��}�(hvK8j  ]�hxh|j  KubK j   )��}�(hvK8j  ]�hxh|j  K ubK!j   )��}�(hvK8j  ]�hxh|j  K!ubK"j   )��}�(hvK8j  ]�hxh|j  K"ubK#j   )��}�(hvK8j  ]�hxh|j  K#ubK$j   )��}�(hvK8j  ]�hxh|j  K$ubK%j   )��}�(hvK8j  ]�hxh|j  K%ubK&j   )��}�(hvK8j  ]�hxh|j  K&ubK'j   )��}�(hvK8j  ]�hxh|j  K'ubK(j   )��}�(hvK8j  ]�hxh|j  K(ubK)j   )��}�(hvK8j  ]�hxh|j  K)ubK*j   )��}�(hvK8j  ]�hxh|j  K*ubK+j   )��}�(hvK8j  ]�hxh|j  K+ubK,j   )��}�(hvK8j  ]�hxh|j  K,ubK-j   )��}�(hvK8j  ]�hxh|j  K-ubK.j   )��}�(hvK8j  ]�hxh|j  K.ubK/j   )��}�(hvK8j  ]�hxh|j  K/ubK0j   )��}�(hvK8j  ]�hxh|j  K0ubK1j   )��}�(hvK8j  ]�hxh|j  K1ubK2j   )��}�(hvK8j  ]�hxh|j  K2ubK3j   )��}�(hvK8j  ]�hxh|j  K3ubK4j   )��}�(hvK8j  ]�hxh|j  K4ubK5j   )��}�(hvK8j  ]�hxh|j  K5ubK6j   )��}�(hvK8j  ]�hxh|j  K6ubK7j   )��}�(hvK8j  ]�hxh|j  K7ubK8j   )��}�(hvK8j  ]�hxh|j  K8ubK9j   )��}�(hvK8j  ]�hxh|j  K9ubK:j   )��}�(hvK8j  ]�hxh|j  K:ubK;j   )��}�(hvK8j  ]�hxh|j  K;ubK<j   )��}�(hvK8j  ]�hxh|j  K<ubK=j   )��}�(hvK8j  ]�hxh|j  K=ubK>j   )��}�(hvK8j  ]�hxh|j  K>ubK?j   )��}�(hvK8j  ]�hxh|j  K?ubK@j   )��}�(hvK8j  ]�hxh|j  K@ubKAj   )��}�(hvK8j  ]�hxh|j  KAubKBj   )��}�(hvK8j  ]�hxh|j  KBubKCj   )��}�(hvK8j  ]�hxh|j  KCubuK9}�(K j   )��}�(hvK9j  ]�hxh|j  K ubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubK	j   )��}�(hvK9j  ]�hxh|j  K	ubK
j   )��}�(hvK9j  ]�hxh|j  K
ubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubKj   )��}�(hvK9j  ]�hxh|j  KubK j   )��}�(hvK9j  ]�hxh|j  K ubK!j   )��}�(hvK9j  ]�hxh|j  K!ubK"j   )��}�(hvK9j  ]�hxh|j  K"ubK#j   )��}�(hvK9j  ]�hxh|j  K#ubK$j   )��}�(hvK9j  ]�hxh|j  K$ubK%j   )��}�(hvK9j  ]�hxh|j  K%ubK&j   )��}�(hvK9j  ]�hxh|j  K&ubK'j   )��}�(hvK9j  ]�hxh|j  K'ubK(j   )��}�(hvK9j  ]�hxh|j  K(ubK)j   )��}�(hvK9j  ]�hxh|j  K)ubK*j   )��}�(hvK9j  ]�hxh|j  K*ubK+j   )��}�(hvK9j  ]�hxh|j  K+ubK,j   )��}�(hvK9j  ]�hxh|j  K,ubK-j   )��}�(hvK9j  ]�hxh|j  K-ubK.j   )��}�(hvK9j  ]�hxh|j  K.ubK/j   )��}�(hvK9j  ]�hxh|j  K/ubK0j   )��}�(hvK9j  ]�hxh|j  K0ubK1j   )��}�(hvK9j  ]�hxh|j  K1ubK2j   )��}�(hvK9j  ]�hxh|j  K2ubK3j   )��}�(hvK9j  ]�hxh|j  K3ubK4j   )��}�(hvK9j  ]�hxh|j  K4ubK5j   )��}�(hvK9j  ]�hxh|j  K5ubK6j   )��}�(hvK9j  ]�hxh|j  K6ubK7j   )��}�(hvK9j  ]�hxh|j  K7ubK8j   )��}�(hvK9j  ]�hxh|j  K8ubK9j   )��}�(hvK9j  ]�hxh|j  K9ubK:j   )��}�(hvK9j  ]�hxh|j  K:ubK;j   )��}�(hvK9j  ]�hxh|j  K;ubK<j   )��}�(hvK9j  ]�hxh|j  K<ubK=j   )��}�(hvK9j  ]�hxh|j  K=ubK>j   )��}�(hvK9j  ]�hxh|j  K>ubK?j   )��}�(hvK9j  ]�hxh|j  K?ubK@j   )��}�(hvK9j  ]�hxh|j  K@ubKAj   )��}�(hvK9j  ]�hxh|j  KAubKBj   )��}�(hvK9j  ]�hxh|j  KBubKCj   )��}�(hvK9j  ]�hxh|j  KCubuK:}�(K j   )��}�(hvK:j  ]�hxh|j  K ubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubK	j   )��}�(hvK:j  ]�hxh|j  K	ubK
j   )��}�(hvK:j  ]�hxh|j  K
ubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubKj   )��}�(hvK:j  ]�hxh|j  KubK j   )��}�(hvK:j  ]�hxh|j  K ubK!j   )��}�(hvK:j  ]�hxh|j  K!ubK"j   )��}�(hvK:j  ]�hxh|j  K"ubK#j   )��}�(hvK:j  ]�hxh|j  K#ubK$j   )��}�(hvK:j  ]�hxh|j  K$ubK%j   )��}�(hvK:j  ]�hxh|j  K%ubK&j   )��}�(hvK:j  ]�hxh|j  K&ubK'j   )��}�(hvK:j  ]�hxh|j  K'ubK(j   )��}�(hvK:j  ]�hxh|j  K(ubK)j   )��}�(hvK:j  ]�hxh|j  K)ubK*j   )��}�(hvK:j  ]�hxh|j  K*ubK+j   )��}�(hvK:j  ]�hxh|j  K+ubK,j   )��}�(hvK:j  ]�hxh|j  K,ubK-j   )��}�(hvK:j  ]�hxh|j  K-ubK.j   )��}�(hvK:j  ]�hxh|j  K.ubK/j   )��}�(hvK:j  ]�hxh|j  K/ubK0j   )��}�(hvK:j  ]�hxh|j  K0ubK1j   )��}�(hvK:j  ]�hxh|j  K1ubK2j   )��}�(hvK:j  ]�hxh|j  K2ubK3j   )��}�(hvK:j  ]�hxh|j  K3ubK4j   )��}�(hvK:j  ]�hxh|j  K4ubK5j   )��}�(hvK:j  ]�hxh|j  K5ubK6j   )��}�(hvK:j  ]�hxh|j  K6ubK7j   )��}�(hvK:j  ]�hxh|j  K7ubK8j   )��}�(hvK:j  ]�hxh|j  K8ubK9j   )��}�(hvK:j  ]�hxh|j  K9ubK:j   )��}�(hvK:j  ]�hxh|j  K:ubK;j   )��}�(hvK:j  ]�hxh|j  K;ubK<j   )��}�(hvK:j  ]�hxh|j  K<ubK=j   )��}�(hvK:j  ]�hxh|j  K=ubK>j   )��}�(hvK:j  ]�hxh|j  K>ubK?j   )��}�(hvK:j  ]�hxh|j  K?ubK@j   )��}�(hvK:j  ]�hxh|j  K@ubKAj   )��}�(hvK:j  ]�hxh|j  KAubKBj   )��}�(hvK:j  ]�hxh|j  KBubKCj   )��}�(hvK:j  ]�hxh|j  KCubuK;}�(K j   )��}�(hvK;j  ]�hxh|j  K ubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�Kahxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubK	j   )��}�(hvK;j  ]�hxh|j  K	ubK
j   )��}�(hvK;j  ]�hxh|j  K
ubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubKj   )��}�(hvK;j  ]�hxh|j  KubK j   )��}�(hvK;j  ]�hxh|j  K ubK!j   )��}�(hvK;j  ]�hxh|j  K!ubK"j   )��}�(hvK;j  ]�hxh|j  K"ubK#j   )��}�(hvK;j  ]�hxh|j  K#ubK$j   )��}�(hvK;j  ]�hxh|j  K$ubK%j   )��}�(hvK;j  ]�hxh|j  K%ubK&j   )��}�(hvK;j  ]�hxh|j  K&ubK'j   )��}�(hvK;j  ]�hxh|j  K'ubK(j   )��}�(hvK;j  ]�hxh|j  K(ubK)j   )��}�(hvK;j  ]�hxh|j  K)ubK*j   )��}�(hvK;j  ]�hxh|j  K*ubK+j   )��}�(hvK;j  ]�hxh|j  K+ubK,j   )��}�(hvK;j  ]�hxh|j  K,ubK-j   )��}�(hvK;j  ]�hxh|j  K-ubK.j   )��}�(hvK;j  ]�hxh|j  K.ubK/j   )��}�(hvK;j  ]�hxh|j  K/ubK0j   )��}�(hvK;j  ]�hxh|j  K0ubK1j   )��}�(hvK;j  ]�hxh|j  K1ubK2j   )��}�(hvK;j  ]�hxh|j  K2ubK3j   )��}�(hvK;j  ]�hxh|j  K3ubK4j   )��}�(hvK;j  ]�hxh|j  K4ubK5j   )��}�(hvK;j  ]�hxh|j  K5ubK6j   )��}�(hvK;j  ]�hxh|j  K6ubK7j   )��}�(hvK;j  ]�hxh|j  K7ubK8j   )��}�(hvK;j  ]�hxh|j  K8ubK9j   )��}�(hvK;j  ]�hxh|j  K9ubK:j   )��}�(hvK;j  ]�hxh|j  K:ubK;j   )��}�(hvK;j  ]�hxh|j  K;ubK<j   )��}�(hvK;j  ]�hxh|j  K<ubK=j   )��}�(hvK;j  ]�hxh|j  K=ubK>j   )��}�(hvK;j  ]�hxh|j  K>ubK?j   )��}�(hvK;j  ]�hxh|j  K?ubK@j   )��}�(hvK;j  ]�hxh|j  K@ubKAj   )��}�(hvK;j  ]�hxh|j  KAubKBj   )��}�(hvK;j  ]�hxh|j  KBubKCj   )��}�(hvK;j  ]�hxh|j  KCubuK<}�(K j   )��}�(hvK<j  ]�hxh|j  K ubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubK	j   )��}�(hvK<j  ]�hxh|j  K	ubK
j   )��}�(hvK<j  ]�hxh|j  K
ubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�Kahxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubKj   )��}�(hvK<j  ]�hxh|j  KubK j   )��}�(hvK<j  ]�hxh|j  K ubK!j   )��}�(hvK<j  ]�hxh|j  K!ubK"j   )��}�(hvK<j  ]�hxh|j  K"ubK#j   )��}�(hvK<j  ]�hxh|j  K#ubK$j   )��}�(hvK<j  ]�hxh|j  K$ubK%j   )��}�(hvK<j  ]�hxh|j  K%ubK&j   )��}�(hvK<j  ]�hxh|j  K&ubK'j   )��}�(hvK<j  ]�hxh|j  K'ubK(j   )��}�(hvK<j  ]�hxh|j  K(ubK)j   )��}�(hvK<j  ]�hxh|j  K)ubK*j   )��}�(hvK<j  ]�hxh|j  K*ubK+j   )��}�(hvK<j  ]�hxh|j  K+ubK,j   )��}�(hvK<j  ]�hxh|j  K,ubK-j   )��}�(hvK<j  ]�hxh|j  K-ubK.j   )��}�(hvK<j  ]�hxh|j  K.ubK/j   )��}�(hvK<j  ]�hxh|j  K/ubK0j   )��}�(hvK<j  ]�hxh|j  K0ubK1j   )��}�(hvK<j  ]�hxh|j  K1ubK2j   )��}�(hvK<j  ]�hxh|j  K2ubK3j   )��}�(hvK<j  ]�hxh|j  K3ubK4j   )��}�(hvK<j  ]�hxh|j  K4ubK5j   )��}�(hvK<j  ]�hxh|j  K5ubK6j   )��}�(hvK<j  ]�hxh|j  K6ubK7j   )��}�(hvK<j  ]�hxh|j  K7ubK8j   )��}�(hvK<j  ]�hxh|j  K8ubK9j   )��}�(hvK<j  ]�hxh|j  K9ubK:j   )��}�(hvK<j  ]�hxh|j  K:ubK;j   )��}�(hvK<j  ]�hxh|j  K;ubK<j   )��}�(hvK<j  ]�hxh|j  K<ubK=j   )��}�(hvK<j  ]�hxh|j  K=ubK>j   )��}�(hvK<j  ]�hxh|j  K>ubK?j   )��}�(hvK<j  ]�hxh|j  K?ubK@j   )��}�(hvK<j  ]�hxh|j  K@ubKAj   )��}�(hvK<j  ]�hxh|j  KAubKBj   )��}�(hvK<j  ]�hxh|j  KBubKCj   )��}�(hvK<j  ]�hxh|j  KCubuK=}�(K j   )��}�(hvK=j  ]�hxh|j  K ubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�Kahxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubK	j   )��}�(hvK=j  ]�hxh|j  K	ubK
j   )��}�(hvK=j  ]�hxh|j  K
ubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�Kahxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�Kahxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubKj   )��}�(hvK=j  ]�hxh|j  KubK j   )��}�(hvK=j  ]�hxh|j  K ubK!j   )��}�(hvK=j  ]�hxh|j  K!ubK"j   )��}�(hvK=j  ]�hxh|j  K"ubK#j   )��}�(hvK=j  ]�hxh|j  K#ubK$j   )��}�(hvK=j  ]�hxh|j  K$ubK%j   )��}�(hvK=j  ]�hxh|j  K%ubK&j   )��}�(hvK=j  ]�hxh|j  K&ubK'j   )��}�(hvK=j  ]�hxh|j  K'ubK(j   )��}�(hvK=j  ]�hxh|j  K(ubK)j   )��}�(hvK=j  ]�hxh|j  K)ubK*j   )��}�(hvK=j  ]�hxh|j  K*ubK+j   )��}�(hvK=j  ]�hxh|j  K+ubK,j   )��}�(hvK=j  ]�hxh|j  K,ubK-j   )��}�(hvK=j  ]�hxh|j  K-ubK.j   )��}�(hvK=j  ]�hxh|j  K.ubK/j   )��}�(hvK=j  ]�hxh|j  K/ubK0j   )��}�(hvK=j  ]�hxh|j  K0ubK1j   )��}�(hvK=j  ]�hxh|j  K1ubK2j   )��}�(hvK=j  ]�hxh|j  K2ubK3j   )��}�(hvK=j  ]�hxh|j  K3ubK4j   )��}�(hvK=j  ]�hxh|j  K4ubK5j   )��}�(hvK=j  ]�hxh|j  K5ubK6j   )��}�(hvK=j  ]�hxh|j  K6ubK7j   )��}�(hvK=j  ]�hxh|j  K7ubK8j   )��}�(hvK=j  ]�hxh|j  K8ubK9j   )��}�(hvK=j  ]�hxh|j  K9ubK:j   )��}�(hvK=j  ]�hxh|j  K:ubK;j   )��}�(hvK=j  ]�hxh|j  K;ubK<j   )��}�(hvK=j  ]�hxh|j  K<ubK=j   )��}�(hvK=j  ]�hxh|j  K=ubK>j   )��}�(hvK=j  ]�hxh|j  K>ubK?j   )��}�(hvK=j  ]�hxh|j  K?ubK@j   )��}�(hvK=j  ]�hxh|j  K@ubKAj   )��}�(hvK=j  ]�hxh|j  KAubKBj   )��}�(hvK=j  ]�hxh|j  KBubKCj   )��}�(hvK=j  ]�hxh|j  KCubuK>}�(K j   )��}�(hvK>j  ]�hxh|j  K ubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�Kahxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubK	j   )��}�(hvK>j  ]�hxh|j  K	ubK
j   )��}�(hvK>j  ]�hxh|j  K
ubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�Kahxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubKj   )��}�(hvK>j  ]�hxh|j  KubK j   )��}�(hvK>j  ]�hxh|j  K ubK!j   )��}�(hvK>j  ]�hxh|j  K!ubK"j   )��}�(hvK>j  ]�hxh|j  K"ubK#j   )��}�(hvK>j  ]�hxh|j  K#ubK$j   )��}�(hvK>j  ]�hxh|j  K$ubK%j   )��}�(hvK>j  ]�hxh|j  K%ubK&j   )��}�(hvK>j  ]�hxh|j  K&ubK'j   )��}�(hvK>j  ]�hxh|j  K'ubK(j   )��}�(hvK>j  ]�hxh|j  K(ubK)j   )��}�(hvK>j  ]�hxh|j  K)ubK*j   )��}�(hvK>j  ]�hxh|j  K*ubK+j   )��}�(hvK>j  ]�hxh|j  K+ubK,j   )��}�(hvK>j  ]�hxh|j  K,ubK-j   )��}�(hvK>j  ]�hxh|j  K-ubK.j   )��}�(hvK>j  ]�hxh|j  K.ubK/j   )��}�(hvK>j  ]�hxh|j  K/ubK0j   )��}�(hvK>j  ]�hxh|j  K0ubK1j   )��}�(hvK>j  ]�hxh|j  K1ubK2j   )��}�(hvK>j  ]�hxh|j  K2ubK3j   )��}�(hvK>j  ]�hxh|j  K3ubK4j   )��}�(hvK>j  ]�hxh|j  K4ubK5j   )��}�(hvK>j  ]�hxh|j  K5ubK6j   )��}�(hvK>j  ]�hxh|j  K6ubK7j   )��}�(hvK>j  ]�hxh|j  K7ubK8j   )��}�(hvK>j  ]�hxh|j  K8ubK9j   )��}�(hvK>j  ]�hxh|j  K9ubK:j   )��}�(hvK>j  ]�hxh|j  K:ubK;j   )��}�(hvK>j  ]�hxh|j  K;ubK<j   )��}�(hvK>j  ]�hxh|j  K<ubK=j   )��}�(hvK>j  ]�hxh|j  K=ubK>j   )��}�(hvK>j  ]�hxh|j  K>ubK?j   )��}�(hvK>j  ]�hxh|j  K?ubK@j   )��}�(hvK>j  ]�hxh|j  K@ubKAj   )��}�(hvK>j  ]�hxh|j  KAubKBj   )��}�(hvK>j  ]�hxh|j  KBubKCj   )��}�(hvK>j  ]�hxh|j  KCubuK?}�(K j   )��}�(hvK?j  ]�hxh|j  K ubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubK	j   )��}�(hvK?j  ]�hxh|j  K	ubK
j   )��}�(hvK?j  ]�hxh|j  K
ubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�Kahxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubKj   )��}�(hvK?j  ]�hxh|j  KubK j   )��}�(hvK?j  ]�hxh|j  K ubK!j   )��}�(hvK?j  ]�hxh|j  K!ubK"j   )��}�(hvK?j  ]�hxh|j  K"ubK#j   )��}�(hvK?j  ]�hxh|j  K#ubK$j   )��}�(hvK?j  ]�hxh|j  K$ubK%j   )��}�(hvK?j  ]�hxh|j  K%ubK&j   )��}�(hvK?j  ]�hxh|j  K&ubK'j   )��}�(hvK?j  ]�Kahxh|j  K'ubK(j   )��}�(hvK?j  ]�hxh|j  K(ubK)j   )��}�(hvK?j  ]�hxh|j  K)ubK*j   )��}�(hvK?j  ]�hxh|j  K*ubK+j   )��}�(hvK?j  ]�hxh|j  K+ubK,j   )��}�(hvK?j  ]�hxh|j  K,ubK-j   )��}�(hvK?j  ]�hxh|j  K-ubK.j   )��}�(hvK?j  ]�hxh|j  K.ubK/j   )��}�(hvK?j  ]�hxh|j  K/ubK0j   )��}�(hvK?j  ]�hxh|j  K0ubK1j   )��}�(hvK?j  ]�hxh|j  K1ubK2j   )��}�(hvK?j  ]�hxh|j  K2ubK3j   )��}�(hvK?j  ]�hxh|j  K3ubK4j   )��}�(hvK?j  ]�hxh|j  K4ubK5j   )��}�(hvK?j  ]�hxh|j  K5ubK6j   )��}�(hvK?j  ]�hxh|j  K6ubK7j   )��}�(hvK?j  ]�hxh|j  K7ubK8j   )��}�(hvK?j  ]�hxh|j  K8ubK9j   )��}�(hvK?j  ]�hxh|j  K9ubK:j   )��}�(hvK?j  ]�hxh|j  K:ubK;j   )��}�(hvK?j  ]�hxh|j  K;ubK<j   )��}�(hvK?j  ]�hxh|j  K<ubK=j   )��}�(hvK?j  ]�hxh|j  K=ubK>j   )��}�(hvK?j  ]�hxh|j  K>ubK?j   )��}�(hvK?j  ]�hxh|j  K?ubK@j   )��}�(hvK?j  ]�hxh|j  K@ubKAj   )��}�(hvK?j  ]�hxh|j  KAubKBj   )��}�(hvK?j  ]�hxh|j  KBubKCj   )��}�(hvK?j  ]�hxh|j  KCubuK@}�(K j   )��}�(hvK@j  ]�hxh|j  K ubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubK	j   )��}�(hvK@j  ]�hxh|j  K	ubK
j   )��}�(hvK@j  ]�hxh|j  K
ubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubKj   )��}�(hvK@j  ]�hxh|j  KubK j   )��}�(hvK@j  ]�hxh|j  K ubK!j   )��}�(hvK@j  ]�hxh|j  K!ubK"j   )��}�(hvK@j  ]�hxh|j  K"ubK#j   )��}�(hvK@j  ]�hxh|j  K#ubK$j   )��}�(hvK@j  ]�Kahxh|j  K$ubK%j   )��}�(hvK@j  ]�Kahxh|j  K%ubK&j   )��}�(hvK@j  ]�hxh|j  K&ubK'j   )��}�(hvK@j  ]�hxh|j  K'ubK(j   )��}�(hvK@j  ]�hxh|j  K(ubK)j   )��}�(hvK@j  ]�hxh|j  K)ubK*j   )��}�(hvK@j  ]�hxh|j  K*ubK+j   )��}�(hvK@j  ]�hxh|j  K+ubK,j   )��}�(hvK@j  ]�hxh|j  K,ubK-j   )��}�(hvK@j  ]�hxh|j  K-ubK.j   )��}�(hvK@j  ]�hxh|j  K.ubK/j   )��}�(hvK@j  ]�hxh|j  K/ubK0j   )��}�(hvK@j  ]�hxh|j  K0ubK1j   )��}�(hvK@j  ]�hxh|j  K1ubK2j   )��}�(hvK@j  ]�hxh|j  K2ubK3j   )��}�(hvK@j  ]�hxh|j  K3ubK4j   )��}�(hvK@j  ]�hxh|j  K4ubK5j   )��}�(hvK@j  ]�hxh|j  K5ubK6j   )��}�(hvK@j  ]�hxh|j  K6ubK7j   )��}�(hvK@j  ]�hxh|j  K7ubK8j   )��}�(hvK@j  ]�hxh|j  K8ubK9j   )��}�(hvK@j  ]�hxh|j  K9ubK:j   )��}�(hvK@j  ]�hxh|j  K:ubK;j   )��}�(hvK@j  ]�hxh|j  K;ubK<j   )��}�(hvK@j  ]�hxh|j  K<ubK=j   )��}�(hvK@j  ]�hxh|j  K=ubK>j   )��}�(hvK@j  ]�hxh|j  K>ubK?j   )��}�(hvK@j  ]�hxh|j  K?ubK@j   )��}�(hvK@j  ]�hxh|j  K@ubKAj   )��}�(hvK@j  ]�hxh|j  KAubKBj   )��}�(hvK@j  ]�hxh|j  KBubKCj   )��}�(hvK@j  ]�hxh|j  KCubuKA}�(K j   )��}�(hvKAj  ]�hxh|j  K ubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubK	j   )��}�(hvKAj  ]�hxh|j  K	ubK
j   )��}�(hvKAj  ]�hxh|j  K
ubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubKj   )��}�(hvKAj  ]�hxh|j  KubK j   )��}�(hvKAj  ]�hxh|j  K ubK!j   )��}�(hvKAj  ]�hxh|j  K!ubK"j   )��}�(hvKAj  ]�Kahxh|j  K"ubK#j   )��}�(hvKAj  ]�hxh|j  K#ubK$j   )��}�(hvKAj  ]�hxh|j  K$ubK%j   )��}�(hvKAj  ]�hxh|j  K%ubK&j   )��}�(hvKAj  ]�hxh|j  K&ubK'j   )��}�(hvKAj  ]�hxh|j  K'ubK(j   )��}�(hvKAj  ]�hxh|j  K(ubK)j   )��}�(hvKAj  ]�hxh|j  K)ubK*j   )��}�(hvKAj  ]�hxh|j  K*ubK+j   )��}�(hvKAj  ]�hxh|j  K+ubK,j   )��}�(hvKAj  ]�hxh|j  K,ubK-j   )��}�(hvKAj  ]�hxh|j  K-ubK.j   )��}�(hvKAj  ]�hxh|j  K.ubK/j   )��}�(hvKAj  ]�hxh|j  K/ubK0j   )��}�(hvKAj  ]�hxh|j  K0ubK1j   )��}�(hvKAj  ]�hxh|j  K1ubK2j   )��}�(hvKAj  ]�hxh|j  K2ubK3j   )��}�(hvKAj  ]�hxh|j  K3ubK4j   )��}�(hvKAj  ]�hxh|j  K4ubK5j   )��}�(hvKAj  ]�hxh|j  K5ubK6j   )��}�(hvKAj  ]�hxh|j  K6ubK7j   )��}�(hvKAj  ]�hxh|j  K7ubK8j   )��}�(hvKAj  ]�hxh|j  K8ubK9j   )��}�(hvKAj  ]�hxh|j  K9ubK:j   )��}�(hvKAj  ]�hxh|j  K:ubK;j   )��}�(hvKAj  ]�hxh|j  K;ubK<j   )��}�(hvKAj  ]�hxh|j  K<ubK=j   )��}�(hvKAj  ]�hxh|j  K=ubK>j   )��}�(hvKAj  ]�hxh|j  K>ubK?j   )��}�(hvKAj  ]�hxh|j  K?ubK@j   )��}�(hvKAj  ]�hxh|j  K@ubKAj   )��}�(hvKAj  ]�hxh|j  KAubKBj   )��}�(hvKAj  ]�hxh|j  KBubKCj   )��}�(hvKAj  ]�hxh|j  KCubuKB}�(K j   )��}�(hvKBj  ]�hxh|j  K ubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubK	j   )��}�(hvKBj  ]�hxh|j  K	ubK
j   )��}�(hvKBj  ]�hxh|j  K
ubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubKj   )��}�(hvKBj  ]�hxh|j  KubK j   )��}�(hvKBj  ]�hxh|j  K ubK!j   )��}�(hvKBj  ]�hxh|j  K!ubK"j   )��}�(hvKBj  ]�hxh|j  K"ubK#j   )��}�(hvKBj  ]�hxh|j  K#ubK$j   )��}�(hvKBj  ]�hxh|j  K$ubK%j   )��}�(hvKBj  ]�hxh|j  K%ubK&j   )��}�(hvKBj  ]�hxh|j  K&ubK'j   )��}�(hvKBj  ]�hxh|j  K'ubK(j   )��}�(hvKBj  ]�hxh|j  K(ubK)j   )��}�(hvKBj  ]�hxh|j  K)ubK*j   )��}�(hvKBj  ]�hxh|j  K*ubK+j   )��}�(hvKBj  ]�hxh|j  K+ubK,j   )��}�(hvKBj  ]�hxh|j  K,ubK-j   )��}�(hvKBj  ]�hxh|j  K-ubK.j   )��}�(hvKBj  ]�hxh|j  K.ubK/j   )��}�(hvKBj  ]�hxh|j  K/ubK0j   )��}�(hvKBj  ]�hxh|j  K0ubK1j   )��}�(hvKBj  ]�hxh|j  K1ubK2j   )��}�(hvKBj  ]�hxh|j  K2ubK3j   )��}�(hvKBj  ]�hxh|j  K3ubK4j   )��}�(hvKBj  ]�hxh|j  K4ubK5j   )��}�(hvKBj  ]�hxh|j  K5ubK6j   )��}�(hvKBj  ]�hxh|j  K6ubK7j   )��}�(hvKBj  ]�hxh|j  K7ubK8j   )��}�(hvKBj  ]�hxh|j  K8ubK9j   )��}�(hvKBj  ]�hxh|j  K9ubK:j   )��}�(hvKBj  ]�hxh|j  K:ubK;j   )��}�(hvKBj  ]�hxh|j  K;ubK<j   )��}�(hvKBj  ]�hxh|j  K<ubK=j   )��}�(hvKBj  ]�hxh|j  K=ubK>j   )��}�(hvKBj  ]�hxh|j  K>ubK?j   )��}�(hvKBj  ]�hxh|j  K?ubK@j   )��}�(hvKBj  ]�hxh|j  K@ubKAj   )��}�(hvKBj  ]�hxh|j  KAubKBj   )��}�(hvKBj  ]�hxh|j  KBubKCj   )��}�(hvKBj  ]�hxh|j  KCubuKC}�(K j   )��}�(hvKCj  ]�hxh|j  K ubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubK	j   )��}�(hvKCj  ]�hxh|j  K	ubK
j   )��}�(hvKCj  ]�hxh|j  K
ubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubKj   )��}�(hvKCj  ]�hxh|j  KubK j   )��}�(hvKCj  ]�hxh|j  K ubK!j   )��}�(hvKCj  ]�hxh|j  K!ubK"j   )��}�(hvKCj  ]�hxh|j  K"ubK#j   )��}�(hvKCj  ]�hxh|j  K#ubK$j   )��}�(hvKCj  ]�hxh|j  K$ubK%j   )��}�(hvKCj  ]�hxh|j  K%ubK&j   )��}�(hvKCj  ]�hxh|j  K&ubK'j   )��}�(hvKCj  ]�hxh|j  K'ubK(j   )��}�(hvKCj  ]�hxh|j  K(ubK)j   )��}�(hvKCj  ]�hxh|j  K)ubK*j   )��}�(hvKCj  ]�hxh|j  K*ubK+j   )��}�(hvKCj  ]�hxh|j  K+ubK,j   )��}�(hvKCj  ]�hxh|j  K,ubK-j   )��}�(hvKCj  ]�hxh|j  K-ubK.j   )��}�(hvKCj  ]�hxh|j  K.ubK/j   )��}�(hvKCj  ]�hxh|j  K/ubK0j   )��}�(hvKCj  ]�hxh|j  K0ubK1j   )��}�(hvKCj  ]�hxh|j  K1ubK2j   )��}�(hvKCj  ]�hxh|j  K2ubK3j   )��}�(hvKCj  ]�hxh|j  K3ubK4j   )��}�(hvKCj  ]�hxh|j  K4ubK5j   )��}�(hvKCj  ]�hxh|j  K5ubK6j   )��}�(hvKCj  ]�hxh|j  K6ubK7j   )��}�(hvKCj  ]�hxh|j  K7ubK8j   )��}�(hvKCj  ]�hxh|j  K8ubK9j   )��}�(hvKCj  ]�hxh|j  K9ubK:j   )��}�(hvKCj  ]�hxh|j  K:ubK;j   )��}�(hvKCj  ]�hxh|j  K;ubK<j   )��}�(hvKCj  ]�hxh|j  K<ubK=j   )��}�(hvKCj  ]�hxh|j  K=ubK>j   )��}�(hvKCj  ]�hxh|j  K>ubK?j   )��}�(hvKCj  ]�hxh|j  K?ubK@j   )��}�(hvKCj  ]�hxh|j  K@ubKAj   )��}�(hvKCj  ]�hxh|j  KAubKBj   )��}�(hvKCj  ]�hxh|j  KBubKCj   )��}�(hvKCj  ]�hxh|j  KCubuu�	tilesSeen�]��djikstra_Stairs_Down�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NKaK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKGKFKEKFKEKDKEKFKGKHKIKJKKKLKMKNKOKPKQKRKSKTKSKTKUKVKWKXKYKZK[K\K]K^K_K`KaKbNe]�(NK`K_K^K]NNKZKYKXKWKVKUKTKSKRKQKPKOKNNKLKKKJKIKHKGKFKEKFKEKDKEKDKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQKRKSKRKSKTKUKVKWKXNKZK[K\K]K^NK`KaNe]�(NK_K^K]K\K[NKYKXKWKVKUNNKRNKPKOKNKMKLKKNKIKHKGKFKEKDKEKDKCKDKCKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQKRKQKRKSKTKUKVKWKXKYKZK[K\K]K^K_K`Ne]�(NK^K]K\NKZKYKXKWNKUKTKSKRKQNKOKNKMKLKKKJKIKHKGKFKEKDKCKDKCKBKCKBKAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQKPKQKRKSKTKUKVKWKXKYKZK[K\K]K^K_Ne]�(NK]K\K[NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKCKBKAKBKAK@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKONKOKPNKTKSKTKUKVKWKXKYNK[K\K]K^Ne]�(NK\K[KZKYKXKWKVKUKTKSKRKQKPNKNKMKLKKKJKIKHKGKFKEKDKCKBKAKBKAK@KAK@K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNNKNKOKPNKRKSKTKUKVKWKXKYKZNK\K]Ne]�(NK[KZKYKXKWKVKUKTKSKRNKPKOKNKMKLKKNKINKGKFKEKDKCKBKAK@KAK@K?K@K?K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMNKMKNKOKPKQKRKSKTKUKVKWKXKYKZK[K\Ne]�(NKZKYNKWKVKUKTKSKRKQKPKONKMKLNKJKIKHKGKFKEKDKCKBKAK@K?K@K?K>K?K>K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKKKLKMNKOKPNKRKSKTKUKVKWKXKYKZK[Ne]�(NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKHNKDKCNNK@K?K>K?K>K=K>K=K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKJKKKLKMKNKONKQKRKSKTKUKVNKXKYKZNe]�(NKXKWKVKUKTKUKTNKPKOKNKMKLNKJKIKHKGKFNKDNKBKAK@K?K>K=NK=K<K=K<K;K<K=K>K?K@KAKBKCNKGKFKGKHKIKJKIKJKKKLKMKNKOKPKQKRNKTKUKVKWKXKYNe]�(NKWKVNKTKSKTNKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@NK>K=K<K=K<K;NNK:K;K<K=K>K?K@KAKBKCNKEKFKGKHKIKHKIKJKKKLKMKNKOKPNKRKSKTKUKVKWKXNe]�(NKVKUKTKSKRNKPKOKNKMKLKMNKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K<K;K:K9K:K9K:K;K<K=K>K?K@KAKBKCKDKEKFKGKHKGKHKIKJKKKLKMKNKOKPKQKRNKTKUKVKWNe]�(NKUKTKSKRKQKPKOKNNKLKKNKINKGKFKEKDKCKBKAK@NK>K=K<K;K:K;K:K9K8NK8K9K:K;K<K=K>K?K@KAKBKCKDNNKGKFKGKHKIKJKKKLKMKNKOKPKQKRKSKTKUKVNe]�(NKTKSKRKQKPKOKNKMKLKKKJNKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK9K8K7K8K7K8K9K:K;K<K=K>K?K@KANKCKDKEKFKEKFKGKHKIKJKKKLKMKNKOKPKQKRKSKTKUNe]�(NKSKRKQKPKOKNKMKLKKKJKIKHKGNKEKDKCKBKANK?K>K=K<K;K:K9K8NNK7K6NK6K7K8K9K:K;K<K=K>K?K@KAKBKCNKEKDKEKFKGKHKIKJKKNKOKNKOKPKQKRKSKTNe]�(NKRKQKPKOKNNKNNKJKIKHKGKFKEKDKCKBKAK@K?NK=K<K;NK9K8K7K6K7K6K5K6K5K6K7K8K9K:K;K<K=K>NK@KAKBKCKDKCKDKEKFKGKHKIKJNKNKMKNKOKPKQKRKSNe]�(NKQKPNKNKMKLKMKLKKKJNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K6K5K4K5K4K5K6K7K8K9K:K;K<K=K>K?K@KAKBNKBKCKDKEKFKGKHKIKJNKLKMKNKOKPKQKRNe]�(NKPKOKNKMKLKKKLKMKLKKNKEKDKCKBKCNK?K>K=K<K;NK9NK7NK5K4K5K4K3K4K3K4K5K6K7K8K9K:K;K<K=K>K?K@KAKBKAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQNe]�(NKOKNKMKLKKKJKKKLNNKENKCKBKANK?K>K=K<K;K:NK8K7K6K5NK3K4K3K2K3K2K3K4K5K6K7K8K9K:K;K<K=K>K?K@KAK@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPNe]�(NKNKMKLKKKJKINNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K3K2K1K2K1K2K3K4K5K6K7K8K9K:K;K<K=K>K?K@K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKONe]�(NKMKLKKNKIKHKGKFKENKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K2K1K0K1K0K1K2K3K4K5K6K7K8K9K:K;K<K=K>K?K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNNe]�(NKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0NK0K/NK/K0K1K2K3K4K5K6K7K8K9K:K;K<K=K>K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMNe]�(NKKKJKIKHNKFKENKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4K3NK1K0K/NK/K.K-K.K/K0K1K2K3K4K5K6K7K8K9K:K;K<K=K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLNe]�(NKJNKHKGKFNKDKCKBKCNK?K>K=K<K;K:K9K8NK6K5K4K3K2K1K0K/K.K/K.K-K,K-K.K/K0K1K2K3K4K5K6K7K8K9K:K;K<K;K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKNe]�(NKIKHKGKFKEKDKCKBKANK?K>K=K<K;K:K9K8K7NK5K4K3K2NK0K/NK-K.K-K,K+K,K-K.K/K0K1K2K3K4K5K6K7K8K9K:K;K:K;K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJNe]�(NKHKGKFKEKDKCKBKAK@K?NK=NNK:K9K8K7K6K5K4K3NK1K0K/K.K-K,K-K,K+K*NNNNNNNNNNNNNNNNK9K:K;K<K=K>K?K@NKDKCKDNKFKGKHKINe]�(NKGKFKEKDKCNKAK@K?K>K=K<K;K:K9K8NK6K5K4K3K2NK0K/K.K-K,K+K,K+K*K)NK+K,K-K.K/K0K1K2K3K4K5K6K7K8NK8K9K:K;K<K=K>K?K@NKBKCKDKEKFKGKHNe]�(NKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K1NK/K.K-K,K+K*K+K*K)K(NK*K+K,K-K.K/K0K1K2K3K4K5K6K7NK7K8K9K:K;K<K=K>K?K@KAKBKCKDKEKFKGNe]�(NKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7NK5K4K3K2K1K0K/K.K-K,K+K*K)K*K)K(K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6NK6K7K8K9K:K;K<K=K>K?K@KAKBKCKDKEKFNe]�(NKDKCKBKAK@NNNK<K;K:NK8NK6K5NK3K2K1K0K/K.K-K,K+K*K)K(K)K(K'K&NK*K+K,K-K.K/K0K1K2K3K4K5K6K7NK5K6K7K8K9K:K;K<NK>K?K@KAKBKCKDKENe]�(NKCKBKAK@K?K>NK<K;K:K9K8K7K6K5K4K3K2NK0K/K.K-K,K+K*K)K(K'K(K'K&K%NK+K,K-K.K/K0K1K2K3K4K5K6K7K8NK4K5K6K7K8K9K:K;K<K=K>K?K@KAKBKCKDNe]�(NKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-NK+K*K)K(K'K&K'K&K%K$NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NK3K4K5K6K7K8K9K:K;K<K=K>K?K@NKDKCNe]�(NKANK?K>NK<K;K:NK8K7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K&K%K$K#NNNNNNNNNNNNNNNNK2K3K4K5K6K7K8K9NK;K<K=K>NK@NKBNe]�(NK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K%NK#K"K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1NNK4K5K6K7K8NK:K;K<K=K>K?K@KANe]�(NK?NK=NK;K:K9K8K7NK5K4K3K2K1NK/K.K-K,K+K*K)K(K'NK%NK#NK#K"K!K K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4NK6K7NK9K:K;K<K=K>K?K@Ne]�(NK>K=K<K;K:NK8K7K6NK4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K#K"K!K KK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6NK8K9K:K;K<NK>K?Ne]�(NK=NNK:K9NK7K6K5K4K3NK1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K"K!K KKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2NK4K5K6K7K8K9K:K;K<K=K>Ne]�(NK<K;K:NK8K7K6K5K4K3K2K1K0K/K.K-K,NNK+NK'K&K%K$K#K"K!K K!K NKKKKK K!K"K#K$K%K&K'K(K)K*K+K,NK.K/K0K1K2K3K4NK6K7NNK:K;K<K=Ne]�(NK;K:K9K8K7K6K5K4K3K2K1K0K/K.NK,K+K*K)NNK&K%K$K#K"K!K KK KKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2NK4K5K6K7K8K9K:K;K<Ne]�(NK:K9K8K7K6K5K4K3K2NK0K/K.K-K,K+NK)K(K'K&K%NK#K"K!K KKNKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+NK-K.K/K0K1K2K3K4K5K6K7K8K9K:K;Ne]�(NK9K8K7K6K5NK3K2K1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!K NKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*NK,K-K.K/K0K1K2K3K4NK6K7K8K9K:Ne]�(NK8K7NK5K4K3K2K1K0K/K.K-K,NK*K)NK'K&K%K$K#K"K!K KKKKKKKNKKKKKNKNK!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7K8K9Ne]�(NK7K6K5K4K3K2NK0NK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKNKKK K!K"K#NK%K&NK(K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7K8Ne]�(NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K"NKKKNKKKKKKKKKKKKKNK K!K"K#K$K%K&K'K(NK*K+K,K-NK/K0K1K2K3K4K5K6K7Ne]�(NK5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$NK"K!K NKKKKKNKKKKKNNKNKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6Ne]�(NK4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#NK!K KNKKKKKKKNKKKKKKKNKKKKKK K!K"NK$K%K&K'K(NK*K+NK-K.K/K0K1K2K3K4K5Ne]�(NK3K2K1K0K/K.K-K,NK*K)K(K'NNNNK"K!K KKKKNKKKKKKKKKKKKKNKKKKKKK K!K"K#K$NK(K'K(K)K*K+K,K-K.K/K0K1K2K3K4Ne]�(NK2K1K0K/K.K-NK+NK)K(K'K&K%K$K#K"K!K KNKKKKNKKKNKKKKKKKKKKKKKKNKK K!NK#K$NK&K'K(NK*K+K,K-K.K/K0K1K2K3Ne]�(NK1K0K/K.NK,NK*K)K(K'K&K%K$K#K"K!K NKKKKKKKKKKNKKKKKKKKKKKKNKKKKK K!K"K#K$K%K&K'NK)K*K+K,K-K.K/K0K1K2Ne]�(NK0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKNKKKNKKKKKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1Ne]�(NK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKNKKKKKKKKKKKKKKKKNKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0Ne]�(NK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKNKKKKKKKKKKKKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/Ne]�(NK-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.Ne]�(NK,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKNKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-Ne]�(NK+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKNKKNKKKKKKKKKKKKKNKKNKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,Ne]�(NK*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKNKKKKKKKKKNKKKNKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+Ne]�(NK)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	K
KKKKKKKKKKKNKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*Ne]�(NK(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KNNNNNNNNKKKKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)Ne]�(NK'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKNK	K
KKKKNKKKKKKKKNKKNKKKKK K!K"K#K$K%K&K'K(Ne]�(NK&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKNKK	K
KKKNKKKKKKKKKKKNKKKKKK K!K"K#K$K%K&K'Ne]�(NK%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKKK	K
KKNKKKKKKKKKKKKNKKNKKK K!K"K#K$K%K&Ne]�(NK$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKNKK	K
KKKNKKKKKKKKNKKKKKKKKKKK K!K"K#K$K%Ne]�(NK#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKNK	K
KKKKNKKKKKKKKKKKKKNKKKKKKK K!K"K#K$Ne]�(NK"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKKNK
KKKKKNKKKKKKKKKKNKKKKKKKKKKK K!K"K#Ne]�(NK!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKKKK NNNNNNNK
KKKKKKKKKKKKKKKKKKKKKK K!K"Ne]�(NK"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKKKKKKKKKKK	K
KKKKKKKKKKKKKKKKKKKKKK K!Ne]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�	eliteList�]��Enemies.Goblins��Goblin_Stonewall���a�
messageSys��
MessageSys��Messages���)��}�(�messages�]�(�Player Ready: Kyle��
Game Start�e�retrieveLimit�K�messageLimit�M�ub�healingList�]�hSa�CollisionMap�]�(]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K KKK K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K KK K Ke]�(KK K K K K KK K K K K KKK KK K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K KK K K K KK K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K KK K K K Ke]�(KK K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K KK K K K K K K K K KK K Ke]�(KK K K K K K K K K K KK K K K K K KK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K Ke]�(KK K KK K K K K K K K K KK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K KK K KKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K Ke]�(KK K K K K K K KK K K K K KK K K K K KK KK K K K K K KK K K K K K K K K K K K K KK K K K K K K K K K K K K K K K KK K K K K K Ke]�(KK K KK K K KK K K K K K K K K K K K K K K K K KK K K K K K KKK K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K Ke]�(KK K K K K KK K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K Ke]�(KK K K K K K K K KK K KK KK K K K K K K K KK K K K K K K K K KK K K K K K K K K K K K K KKK K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K KK K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K KK K K K K KK K K K K K K K KKK K KK K K K K K K K K K K K K K KK K K K K K K K K KK K K K K K K K Ke]�(KK K K K K KK KK K K K K K K K K K K K KK K K KK K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K KK K K K K K K K Ke]�(KK K KK K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K KK K K K K K K Ke]�(KK K K K K K K K K K KK K K K K KK K K K K KK KK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K KKK KK K K KK K K K K K KK K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K KKK K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K KK K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K KK K KK K K K K K K K K K K KK K K K K KK K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK KK K K KK K K K KK K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K KK K K K K K K K K KK K K K KK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K KK KKK K K K K K K K KK K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K KK K K KK K K K Ke]�(KK K K K K KK K K K K K K K K K KK K K K K KK K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K KK K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K KK K K K KK K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K Ke]�(KK K K K K KKKK K K KK KK K KK K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K KK K K K K K K K Ke]�(KK K K K K K KK K K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K KK K Ke]�(KK KK K KK K K KK K K K K K K K K K K K K K KK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K KK K K K KK KK Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K KKK K K K K KK K K K K K K K Ke]�(KK KK KK K K K K KK K K K K KK K K K K K K K K KK KK KK K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K Ke]�(KK K K K K KK K K KK K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K KK K Ke]�(KK KKK K KK K K K K KK K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K Ke]�(KK K K KK K K K K K K K K K K K K KKK KK K K K K K K K K K KK K K K K K K K K K K K K K K K K KK K K K K K K KK K KKK K K K Ke]�(KK K K K K K K K K K K K K K KK K K K KKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K Ke]�(KK K K K K K K K K KK K K K K K KK K K K K KK K K K K K KK K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K Ke]�(KK K K K K KK K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K KK K K K K Ke]�(KK K KK K K K K K K K K K KK K KK K K K K K K K K K K K K K K KK K K K K KK KK K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K KK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K KK K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K KK K K K K K KK K K KK K K K K K K K K K K K K KK K K K K K K K K KK K K K KK K K K K K K K K Ke]�(KK K K K K K K K K K K K K K KK K K KK K K KK K K K K KK K K K K KKK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K KK K K KK K K K K K K KK K K K K K K KK K K K K K K K KK K K K K KK K KK K K K K K K K K Ke]�(KK K K K K K K K KK K K K KKKKK K K K K K K KK K K K K K K K K K K K K KK K K K K K K K K K K KK K K K K K K K K K K K K K K Ke]�(KK K K K K K KK KK K K K K K K K K K K KK K K K KK K K KK K K K K K K K K K K K K K KK K K KK K KK K K KK K K K K K K K K K Ke]�(KK K K K KK KK K K K K K K K K K K KK K K K K K K K K K KK K K K K K K K K K K K KK K K K K K K K K K K K KK K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K K K K K K KK K KK K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K KK K K KK K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K KK K KK K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K K K K KK K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K KK K KK K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K KK K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K K K K K K KK K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K K K KK K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKee�	enemyList�]�(j�8  �Goblin_Lancer���j�8  �Goblin_Berserker���j�8  �Goblin_Archer���j�8  �Goblin_Knight���j�8  �Goblin_Grunt���j�8  �Goblin_Thief���e�textWall��Bricks
��	equipList�]�(h	h�Iron_Shield���h�Buckler���h�Wooden_Shield���h�	Longsword���h�
Greatsword���h�Bow���h�Spear���h�Dagger���hg�Cloth_Shirt���hihg�Leather_Shirt���hg�Leather_Helm���hg�Iron_Breastplate���hg�	Iron_Helm���hg�Chain_Shirt���hg�
Chain_Helm���ehqht�djikstra_Player�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NK G�\������G�\�     G�\333333G�[�fffffG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�F������G�F333333G�E������G�E      G�DffffffNe]�(NG�\������G�\�     G�\333333G�[�fffffNNG�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffNG�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      NG�F������G�F333333G�E������G�F333333G�E������NG�DffffffG�C������Ne]�(NG�\�     G�\333333G�[�fffffG�[������G�[L�����NG�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     NNG�X������NG�X      G�W�33333G�WffffffG�W�����G�V������G�V�     NG�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S�����͕      G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�E������G�E      G�DffffffG�C������G�C333333Ne]�(NG�\333333G�[�fffffG�[������NG�[      G�Z�33333G�ZffffffG�Z�����NG�Y�     G�Y333333G�X�fffffG�X������G�XL�����NG�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�E      G�DffffffG�C������G�C333333G�B������Ne]�(NG�[�fffffG�[������G�[L�����NG�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      NG�I������G�I333333NG�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������NG�C������G�C333333G�B������G�B      Ne]�(NG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      NG�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffNG�I333333G�H������G�H      NG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�C������G�C333333NG�B      G�AffffffNe]�(NG�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������NG�X      G�W�33333G�WffffffG�W�����G�V������G�V�     NG�U�fffffNG�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������NG�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�C333333G�B������G�B      G�AffffffG�@������Ne]�(NG�[      G�Z�33333NG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333NG�W�����G�V������NG�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffNG�F333333G�E������NG�DffffffG�C������G�C333333G�B������G�B      G�B������G�B      G�AffffffG�@������G�@333333Ne]�(NG�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U������NG�TffffffG�T�����NNG�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      NG�C������G�C333333G�B������G�B      G�AffffffG�B      NG�@������G�@333333G�?333333Ne]�(NG�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�Y�     G�Y333333NG�X      G�W�33333G�WffffffG�W�����G�V������NG�V333333G�U�fffffG�U������G�UL�����G�U      NG�TffffffNG�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����NG�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333NG�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�C333333NG�@������G�AffffffG�@������G�@333333G�?333333G�>      Ne]�(NG�Z�����G�Y������NG�Y333333G�X�fffffG�Y333333NG�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333NG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����NNG�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      NG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      NG�@������G�@333333G�@������G�@333333G�?333333G�>      G�<������Ne]�(NG�Y������G�Y�     G�Y333333G�X�fffffG�X������NG�X      G�W�33333G�WffffffG�W�����G�V������G�W�����NG�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333NG�?333333G�>      G�<������G�;������Ne]�(NG�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffNG�V������G�V�     NG�U�fffffNG�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333NG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333NG�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      NNG�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�?333333G�>      G�<������G�;������G�:ffffffNe]�(NG�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333NG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����NG�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������NG�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�>      G�<������G�;������G�:ffffffG�9333333Ne]�(NG�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����NG�T�33333G�TffffffG�T�����G�S������G�S�     NG�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������NNG�O������G�O333333NG�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333NG�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333NG�>      G�<������G�;������G�<������G�;������G�:ffffffG�9333333G�8      Ne]�(NG�X������G�XL�����G�X      G�W�33333G�WffffffNG�WffffffNG�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffNG�RL�����G�R      G�Q�33333NG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      NG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333NG�<������G�;������G�:ffffffG�;������G�:ffffffG�9333333G�8      G�6������Ne]�(NG�XL�����G�X      NG�WffffffG�W�����G�V������G�W�����G�V������G�V�     G�V333333NG�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffNG�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������NG�:ffffffG�9333333G�:ffffffG�9333333G�8      G�6������G�5������Ne]�(NG�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V������G�W�����G�V������G�V�     NG�T�33333G�TffffffG�T�����G�S������G�T�����NG�R�fffffG�R������G�RL�����G�R      G�Q�33333NG�Q�����NG�P�     NG�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�9333333G�8      G�6������G�5������G�4ffffffNe]�(NG�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�V�     G�V������NNG�T�33333NG�T�����G�S������G�S�     NG�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffNG�P������G�P�     G�P333333G�O������NG�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�8      G�6������G�5������G�4ffffffG�3333333Ne]�(NG�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffNNG�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333NG�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�6������G�5������G�4ffffffG�3333333G�2      Ne]�(NG�W�����G�V������G�V�     NG�U�fffffG�U������G�UL�����G�U      G�T�33333NG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�5������G�4ffffffG�3333333G�2      G�0������Ne]�(NG�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������NG�K������G�K      NG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�4ffffffG�3333333G�2      G�0������G�/333333Ne]�(NG�W�����G�V������G�V�     G�V333333NG�U������G�UL�����NG�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333NG�P�     G�P333333G�O������G�O333333G�N������NG�MffffffG�L������G�L333333NG�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�3333333G�2      G�0������G�/333333G�,������Ne]�(NG�WffffffNG�V������G�V�     G�V333333NG�U������G�UL�����G�U      G�T�33333NG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      NG�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�2      G�0������G�/333333G�,������G�*ffffffNe]�(NG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333NG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333NG�P�     G�P333333G�O������G�O333333NG�N      G�MffffffNG�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�0������G�/333333G�,������G�*ffffffG�(      Ne]�(NG�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����NG�S�     NNG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     NG�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333NNNNNNNNNNNNNNNNG�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333NG�0������G�/333333G�,������NG�,������G�*ffffffG�(      G�%������Ne]�(NG�V�     G�V333333G�U�fffffG�U������G�UL�����NG�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      NG�QffffffG�Q�����G�P������G�P�     G�P333333NG�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������NG�K      G�K������G�L333333G�L������G�MffffffG�N      G�N������G�O333333G�O������G�P333333G�P�     G�P������G�Q�����G�QffffffNG�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������NG�,������G�*ffffffG�(      G�*ffffffG�(      G�%������G�#333333Ne]�(NG�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffNG�P������G�P�     G�P333333G�O������NG�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333NG�JffffffG�K      G�K������G�L333333G�L������G�MffffffG�N      G�N������G�O333333G�O������G�P333333G�P�     G�P������G�Q�����NG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�(      G�%������G�#333333G� ������Ne]�(NG�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����NG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�I333333G�I������G�JffffffG�K      G�K������G�L333333G�L������G�MffffffG�N      G�N������G�O333333G�O������G�P333333G�P�     G�P������NG�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�#333333G�%������G�#333333G� ������G�������Ne]�(NG�V333333G�U�fffffG�U������G�UL�����G�U      NNNG�S������G�S�     G�S333333NG�R������NG�R      G�Q�33333NG�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      NG�JffffffG�K      G�K������G�L333333G�L������G�MffffffG�N      G�N������G�O333333G�O������G�P333333G�P�     G�P������G�Q�����NG�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������NG�(      G�%������G�#333333G� ������G�#333333G� ������G�������G�      Ne]�(NG�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffNG�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������NG�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffNG�K      G�K������G�L333333G�L������G�MffffffG�N      G�N������G�O333333G�O������G�P333333G�P�     G�P������G�Q�����G�QffffffNG�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�#333333G� ������G�������G� ������G�������G�      G�333333Ne]�(NG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������NG�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������NG�K������G�L333333G�L������G�MffffffG�N      G�N������G�O333333G�O������G�P333333G�P�     G�P������G�Q�����G�QffffffG�Q�33333NG�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�#333333G� ������G�������G�      G�������NG�333333G�������Ne]�(NG�UL�����NG�T�33333G�TffffffNG�S������G�S�     G�S333333NG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffNG�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333NNNNNNNNNNNNNNNNG�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffNG� ������G�������G�      G�333333NG�333333NG�333333Ne]�(NG�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������NG�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������NNG�3333333G�2      G�0������G�/333333G�,������NG�������G�      G�333333G�������G�333333G��333333G�       G��333333Ne]�(NG�UL�����NG�T�33333NG�T�����G�S������G�S�     G�S333333G�R�fffffNG�RL�����G�R      G�Q�33333G�QffffffG�Q�����NG�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      NG�I������NG�H������NG�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333NG�0������G�/333333NG� ������G�������G�      G�333333G�������G�333333G��333333G�333333Ne]�(NG�U������G�UL�����G�U      G�T�33333G�TffffffNG�S������G�S�     G�S333333NG�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������NG�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������NG�#333333G� ������G�������G�      G�333333NG�333333G�������Ne]�(NG�U�fffffNNG�TffffffG�T�����NG�S�     G�S333333G�R�fffffG�R������G�RL�����NG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������NG�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333NG�,������G�*ffffffG�(      G�%������G�#333333G� ������G�������G�      G�333333G�������G�333333Ne]�(NG�U������G�UL�����G�U      NG�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333NNG�N������NG�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      NG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffNG�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������NG�(      G�%������NNG�������G�      G�333333G�      Ne]�(NG�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffNG�P������G�P�     G�P333333G�O������NNG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������NG�,������G�*ffffffG�(      G�%������G�#333333G� ������G�������G�      G�������Ne]�(NG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333NG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����NG�O������G�O333333G�N������G�N      G�MffffffNG�L333333G�K������G�K      G�JffffffG�I������G�I333333NG�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333NG�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�#333333G� ������G�������G� ������Ne]�(NG�U�fffffG�U������G�UL�����G�U      G�T�33333NG�T�����G�S������G�S�     G�S333333G�R�fffffNG�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������NG�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffNG�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������NG�(      G�%������G�#333333G� ������G�#333333Ne]�(NG�V333333G�U�fffffNG�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      NG�QffffffG�Q�����NG�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������NG�GffffffG�F������G�F333333G�E������G�E      NG�C������NG�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�#333333G�%������Ne]�(NG�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffNG�S������NG�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������NG�DffffffG�C������G�C333333G�B������G�B      G�AffffffNG�@333333G�?333333NG�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�(      Ne]�(NG�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333NG�Q�����G�P������G�P�     G�P333333G�O������G�O333333NG�N      G�MffffffG�L������NG�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffNG�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������NG�:ffffffG�9333333G�8      G�6������NG�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�*ffffffNe]�(NG�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������NG�R      G�Q�33333G�QffffffNG�P������G�P�     G�P333333NG�O333333G�N������G�N      G�MffffffG�N      NG�K������G�K      G�JffffffG�I������G�I333333NNG�GffffffNG�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�,������Ne]�(NG�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333NG�Q�����G�P������G�P�     NG�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333NG�K      G�JffffffG�I������G�I333333G�H������G�H      G�H������NG�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      NG�@������G�@333333G�?333333G�>      G�<������NG�:ffffffG�9333333NG�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�/333333Ne]�(NG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      NG�TffffffG�T�����G�S������G�S�     NNNNG�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333NG�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�I333333NG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������NG�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�0������Ne]�(NG�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffNG�UL�����NG�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333NG�Q�����G�P������G�P�     G�P������NG�O333333G�N������G�N      NG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      NG�C������G�C333333G�B������NG�AffffffG�B      NG�?333333G�>      G�<������NG�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�2      Ne]�(NG�W�33333G�WffffffG�W�����G�V������NG�V333333NG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������NG�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������NG�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������NG�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      NG�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�3333333Ne]�(NG�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333NG�O333333G�N������G�N      NG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�4ffffffNe]�(NG�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     NG�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������NG�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�5������Ne]�(NG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����NG�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�6������Ne]�(NG�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�8      Ne]�(NG�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333NG�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�9333333Ne]�(NG�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      NG�QffffffG�Q�����NG�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������NG�H������G�H      NG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�:ffffffNe]�(NG�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     NG�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      NG�I������G�I333333G�H������NG�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�;������Ne]�(NG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������NG�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�<������Ne]�(NG�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������NNNNNNNNG�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�>      Ne]�(NG�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����NG�R�fffffG�S333333G�S�     G�S������G�T�����G�TffffffNG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������NG�GffffffG�F������NG�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�?333333Ne]�(NG�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffNG�R������G�R�fffffG�S333333G�S�     G�S������G�T�����NG�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffNG�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�@333333Ne]�(NG�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�R      G�RL�����G�R������G�R�fffffG�S333333G�S�     G�S������NG�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�H������NG�F333333G�E������NG�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�@������Ne]�(NG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      NG�R������G�R�fffffG�S333333G�S�     G�S������G�T�����NG�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffNG�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�AffffffNe]�(NG�[�fffffG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����NG�R�fffffG�S333333G�S�     G�S������G�T�����G�TffffffNG�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      NG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�B      Ne]�(NG�\333333G�[�fffffG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������NG�S333333G�S�     G�S������G�T�����G�TffffffG�T�33333NG�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffNG�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�B������Ne]�(NG�\�     G�\333333G�[�fffffG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�S333333NNNNNNNG�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�C333333Ne]�(NG�\������G�\�     G�\333333G�[�fffffG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�C������Ne]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�levelManager��LevelManager�j�9  ��)��}�(�	gameState��__main__��Game���)��}�(�width�K#�loadRequest���yConst�KK�turn�Kh�h�	levelList�j�9  �MessageHandler�j�8  �height�K�gameVersion��0.1.0��console��tdl��Console���)��KYKE]�(K K K K ��K K K ����KKK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KLK�K�K���K K K ����KEK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KRK�K�K���K K K ����KPK�K�K���K K K ����KAK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KWK�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KGK�K�K���K K K ����KPK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KxK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KaK�K�K���K K K ����KoK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����KFK�K�K���K K K ����K K K K ��K K K ����KvK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KnK�K�K���K K K ����KwK�K�K���K K K ����KmK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KmK�K�K���K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KwK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K0K�K�K���K K K ����K K K K ��K K K ����KhK�K�K���K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K:K�K�K���K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KSK�K�K���K K K ����KrK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KPK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KtK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K1K�K�K���K K K ����K2K�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����KRK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K9K�K�K���K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KrK�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KBK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KtK�K�K���K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KFK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����e(K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KKK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K �����       K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����e(K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����e(K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K@KKYK���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����e(K K�K�K���K K K ����K K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K����       K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����e(K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����e��b�xConst�K,ubj�9  ]�h|aj�8  j�8  �nextSeed�M�M�cursor�K ub�inSeed�M��	textSpace��ground, covered in leaves
��maze�]�(]�(�T�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  �.�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �~�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  hj��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �x�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  hWj��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �#�jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �D�j��  j��  j��  j��  j��  j��  j��  j��  �=�j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  hj��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �X�j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �S�j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  hWj��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jρ  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j́  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  hWj��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jˁ  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jρ  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  hj��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  hWj��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jǁ  j��  jρ  j��  j��  j��  j��  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �E�jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  jǁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  ee�djikstra_Player_Away�jH9  �SeesMap�]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK KK K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K Ke]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK KKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK KKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K KKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKK K K K K KKKK e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K KKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K ee�args�]�(KKe�SeenMap�]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK KK K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K Ke]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK KKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K �2�      K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK KKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K KKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKK K K K K KKKK e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K KKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K eej�9  j�9  �djikstra_Stairs_Up�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NKaK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K&K%K$K#K"Ne]�(NK`K_K^K]NNKZKYKXKWKVKUKTKSKRKQKPKOKNNKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K%K$NK"K!Ne]�(NK_K^K]K\K[NKYKXKWKVKUNNKRNKPKOKNKMKLKKNKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K$K#K"K!K Ne]�(NK^K]K\NKZKYKXKWNKUKTKSKRKQNKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K#K"K!K KNe]�(NK]K\K[NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-NK+K*NK(K'K&K%K$K#K"K!NK!K KKNe]�(NK\K[KZKYKXKWKVKUKTKSKRKQKPNKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,NK*K)K(NK&K%K$K#K"K!K K!K NKKNe]�(NK[KZKYKXKWKVKUKTKSKRNKPKOKNKMKLKKNKINKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K!K KK KKKKNe]�(NKZKYNKWKVKUKTKSKRKQKPKONKMKLNKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$NK"K!K KKKKKKKNe]�(NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKHNKDKCNNK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#NK!K KKKKNKKKNe]�(NKXKWKVKUKTKUKTNKPKOKNKMKLNKJKIKHKGKFNKDNKBKAK@K?K>K=NK;K:K9K8K7K6K5K4K3K2K1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!K KK NKKKKKKNe]�(NKWKVNKTKSKTNKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@NK>K=K<K;K:K9NNK6K5K4K3K2K1K0K/K.K-NK+K*K)K(K'K&K%K$K#K"K!K KKNKKKKKKKNe]�(NKVKUKTKSKRNKPKOKNKMKLKMNKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKNKKKKNe]�(NKUKTKSKRKQKPKOKNNKLKKNKINKGKFKEKDKCKBKAK@NK>K=K<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+K*K)K(NNK%K$K#K"K!K KKKKKKKKKKKKNe]�(NKTKSKRKQKPKOKNKMKLKKKJNKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4K3K2K1K0K/K.K-K,K+K*K)NK'K&K%K$K#K"K!K KKKKKKKKKKKKKNe]�(NKSKRKQKPKOKNKMKLKKKJKIKHKGNKEKDKCKBKANK?K>K=K<K;K:K9K8NNK5K4NK2K1K0K/K.K-K,K+K*K)K(K'K&K%NK#K"K!K KKKKKNKKKKKKKKNe]�(NKRKQKPKOKNNKNNKJKIKHKGKFKEKDKCKBKAK@K?NK=K<K;NK9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K KKKKKKNKKKKKKKKNe]�(NKQKPNKNKMKLKMKLKKKJNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"NK KKKKKKKKNKKKKKKKNe]�(NKPKOKNKMKLKKKLKMKLKKNKEKDKCKBKCNK?K>K=K<K;NK9NK7NK5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKNe]�(NKOKNKMKLKKKJKKKLNNKENKCKBKANK?K>K=K<K;K:NK8K7K6K5NK3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKNe]�(NKNKMKLKKKJKINNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKNe]�(NKMKLKKNKIKHKGKFKENKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKNe]�(NKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0NK.K-NK+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKNe]�(NKMKLKKKJNKHKGNKEKDKCKBKAK@K?K>K=K<K;NK7K6K5K4K3NK1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKNe]�(NKNNKLKKKJNKHKGKFKENKCKBKAK@K?K>K=K<NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKNe]�(NKMKLKKKJKIKHKGKFKENKCKBKAK@K?K>K=K<K;NK7K6K5K4NK2K1NK-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKK
Ne]�(NKLKKKJKIKHKGKFKEKDKCNKANNK>K=K<K;K:K9K8K7NK3K2K1K0K/K.K-K,K+K*NNNNNNNNNNNNNNNNKKKKKKKKNKKKNKKK
K	Ne]�(NKKKJKIKHKGNKEKDKCKBKAK@K?K>K=K<NK:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+NK-K.K/K0K1K2K3K4K5K6K7K8K9K:NKKKKKKKKKNKKK
KK
K	KNe]�(NKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK8K7K6K5NK3K2K1K0K/K.K-K,K+K*NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NKKKKKKKKKKKK
K	K
K	KKNe]�(NKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=NK9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7K8NKKKKKKKKKKK
K	KK	KKKNe]�(NKJKIKHKGKFNNNKBKAK@NK>NK<K;NK7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NKKKKKKKKNK
K	KKKKKKNe]�(NKIKHKGKFKEKDNKBKAK@K?K>K=K<K;K:K9K8NK4K3K2K1K0K/K.K-K,K+K*K)K(K'NK-K.K/K0K1K2K3K4K5K6K7K8K9K:NKKKKKKKKK
K	KKKKKKKNe]�(NKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3NK/K.K-K,K+K*K)K(K'K&NK.K/K0K1K2K3K4K5K6K7K8K9K:K;NKKKKKKKK
K	KKKKKNKKNe]�(NKGNKEKDNKBKAK@NK>K=K<K;K:K9K8K7K6K5K4K3K2K1NK-K,K+K*K)K(K'K&K%NNNNNNNNNNNNNNNNKKKKKKKKNKKKKNKNKNe]�(NKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)NK%K$K#K"K!K KKKKKKKKKKKKKNNKKKKKNKKKKKKK KNe]�(NKGNKENKCKBKAK@K?NK=K<K;K:K9NK5K4K3K2K1K0K/K.K-NK+NK)NK'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKNKKNKKKKKKKKNe]�(NKHKGKFKEKDNKBKAK@NK<K;K:K9K8K7K6K5K4K3NK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKNKKKKKNKKNe]�(NKINNKDKCNKAK@K?K>K=NK9K8K7K6K5K4K3K2K1K0NK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKNKKK
K	KKKKKKKNe]�(NKHKGKFNKBKAK@K?K>K=K<K;K:K9K8K7K6NNK3NK1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K KKKKKKKKKKNKKKKKKKNK
K	NNKKKKNe]�(NKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK8K7K6K5NNK0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKNKKK
K	KKKKKNe]�(NKHKGKFKEKDKCKBKAK@NK>K=K<K;K:K9NK5K4K3K2K1NK/K.K-K,K+K*NK(K'K&K%K$K#K"K!K KKKKKKKKKKKNKKKKKKKKKK
K	KKKKNe]�(NKIKHKGKFKENKCKBKAK@K?NK;K:K9K8K7K6K5K4K3K2K1K0K/K.NK,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKNKKKKKKKKKNK
K	KKKNe]�(NKJKINKEKDKCKBKAK@K?K>K=K<NK:K9NK7K6K5K4K3K2K1K0K/K.K-K,K+K*K)NK'K&K%K$K#NK!NKKKKKKKKKKKKKKKKKKKKKK
K	KK	Ne]�(NKIKHKGKFKEKDNKBNK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$NK"K!K KKKNKKNKKKKKKKKKKKKKKK
K	K
Ne]�(NKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;NK9K8K7K6K5K4NK2K1K0NK.K-K,K+K*K)K(K'K&K%K$K#K"NK KKKKKKKKNKKKKNKKKKKKKK
KNe]�(NKKKJKIKHKGKFKEKDKCKBKAK@K?K>NK<K;K:NK8K7K6NK4K3K2K1K2NK.K-K,K+K*NNK'NK%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKNe]�(NKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;NK9K8K7NK5K4K3K2K1K0K/NK-K,K+K*K)K(K)NK%K$K#K"K!K KKNKKKKKNKKNKKKKKKKKKNe]�(NKMKLKKKJKIKHKGKFNKDKCKBKANNNNK<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+K*K)K*NK&K%K$K#K"K!K KKKKNKKKKKKKKKKKKKKKNe]�(NKNKMKLKKKJKINKGNKEKDKCKBKAK@K?K>K=K<K;NK9K8K7K8NK4K3K2NK0K/K.K-K,K+K*K)K(K'K&K%K$K#NK!K KNKKNKKKNKKKKKKKKKKNe]�(NKOKNKMKLNKJNKHKGKFKEKDKCKBKAK@K?K>NK<K;K:K9K8K7K6K5K4K3NK1K0K/K.K-K,K+K*K)K(K'K&NK$K#K"K!K KKKKKKKNKKKKKKKKKKNe]�(NKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2NK0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKNe]�(NKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7NK5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&NK$K#K"K!K KKKKKKKKKKKKKKKKNe]�(NKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKNe]�(NKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKNe]�(NKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*NK(K'K&K%K$K#K"K!K KKKKKKKKKKKKKNe]�(NKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NK:K9NK7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(NK&K%K$K#K"K!K KKKKKKKKKKKKNe]�(NKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7NK5K4K3K2K1K0K/K.K-NK+K*K)NK'K&K%K$K#K"K!K KKKKKKKKKKKNe]�(NKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K!K KKKKKKKKKKNe]�(NKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8NNNNNNNNK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKNe]�(NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK?K@KAKBKCKDNK0K/K.K-K,K+K*K)NK'K&NK$K#K"K!K KKKKKKKKNe]�(NKZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK>K?K@KAKBKCNK1K0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K KKKKKKKNe]�(NK[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K<K=K>K?K@KAKBNK2K1K0K/K.K-K,K+K*K)K(K)NK%K$NK"K!K KKKKKKNe]�(NK\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NK>K?K@KAKBKCNK3K2K1K0K/K.K-K,NK*K)K(K'K&K%K$K#K"K!K KKKKKNe]�(NK]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=NK?K@KAKBKCKDNK4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K KKKKNe]�(NK^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>NK@KAKBKCKDKENK5K4K3K2K1K0K/K.K-K,NK*K)K(K'K&K%K$K#K"K!K KKKNe]�(NK_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K@NNNNNNNK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KK Ne]�(NK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K K!Ne]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�stairsUp�]�(K"KAe�itemList�]�(hShQ�Bundle_Of_Arrows���hQ�	Time_Bomb���hQ�Scroll_of_Fireball���hQ�Scroll_of_Lightning_Bolt���h	j*9  j,9  j.9  j09  j29  j49  j69  j89  j:9  hij<9  j>9  j@9  jB9  jD9  jF9  ej  }�(K hs)��}�(hvKhwK hhhxh|j  K'h�Item�hrj49  )��}�(hqj؂  hKhKhKhhhhh�h�hKh�hhhKh�hKh�Bow�h�ububKhs)��}�(hvKhwKhj��  hxh|j  K#h�Enemy�hrj9  )��}�(hK
hK hj49  )��}�(hKhKhKhhhhh�h�hKh�hhhKh�hKhj݂  h�ubhKh�h ��isAfraid��h!Kh"�hj��  h-K	hKh.K hK hfhi)��}�(h�h�hKhhhKh.Kh�hhhhlhhmub�	cowardice�G?�      h\KhDN�lastPlayerMap�Nhd]�hFKdhHKh�Goblin Archer�hJK hO]�hCK h]]�h]�(K�KKe�lastPlayerLoc�Nh`K �
dropChance�K(�
stealthVal�K �necklace�NhE�hcNhnKho��hearingDist�Khqjނ  �armor�j<9  )��}�(h�h�hKhhhKh.Kh�hhh�Leather Shirt�h�armor�ub�
alliesList�]�(jނ  hs)��}�(hvKhwKhj��  hxh|j  K'hj��  hrj 9  )��}�(hKhK hj09  )��}�(hKhKhKhhh�1H�h�h�hKh�hhhKh�hKh�	Longsword�h�ubhKh�h �j�  �h!K h"�hj��  h-KhKh.K hK hfjB9  )��}�(h�h�hKhhhKh.Kh�hhh�	Iron Helm�hhmubj�  G        h\KhDNj�  Nhd]�hFKdhHKh�Goblin Knight�hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqj��  j�  j<9  )��}�(h�h�hKhhhKh.Kh�hhhj��  hj��  ubj��  ]�(jނ  j��  e�leftHand�j.9  )��}�(hKhKhhhj�  h�h�h�h�hhhKh.Kh�hK h�Wooden Shield�hK ub�blocking��hKububej�  Nj�  �hKububKj��  Khs)��}�(hvKhwKhj��  hxh|j  K8hj��  hrj"9  )��}�(hK	hK hj09  )��}�(hKhKhKhhhj�  h�h�hKh�hhhKh�hKhj�  h�ubhKh�h �j�  �h!K h"�hj��  h-KhKh.K hK hfj>9  )��}�(h�h�hKhhhKh.K
h�hhh�Leather Helm�hhmubj�  G?��Q�h\KhDNj�  Nhd]�hFKdhHKh�Goblin Grunt�hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqj�  j�  j<9  )��}�(h�h�hKhhhKh.Kh�hhhj��  hj��  ubj��  ]�(j�  hs)��}�(hvKhwKhj��  hxh|j  K6hj��  hrj9  )��}�(hKhK hj29  )��}�(hKhKhKhhhhh�h�hKh�hhhKh�hKh�
Greatsword�h�ubhKh�h �j�  �h!K h"�hj��  h-KhKh.K hK hfj>9  )��}�(h�h�hKhhhKh.K
h�hhhj�  hhmubj�  G        h\KhDNj�  Nhd]�hFKdhHKh�Goblin Berserker�hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqj"�  j�  j<9  )��}�(h�h�hKhhhKh.Kh�hhhj��  hj��  ubj��  ]�(j�  j"�  ej�  Nj�  �hKububej�  Nj�  �hKububKhs)��}�(hvKhwKhhWhxh|j  K5h�Health�hrhS)��}�(hVKh�h�hhWhqj2�  hhhhXhhYububKj"�  Khs)��}�(hvKhwKhj��  hxh|j  K(hj��  hrj9  )��}�(hK
hK hj49  )��}�(hKhKhKhhhhh�h�hKh�hhhKh�hKhj݂  h�ubhKh�h �j�  �h!Kh"�hj��  h-KhKh.K hK hfhi)��}�(h�h�hKhhhKh.Kh�hhhhlhhmubj�  G?�      h\KhDNj�  Nhd]�hFKdhHKhj�  hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqj7�  j�  j<9  )��}�(h�h�hKhhhKh.Kh�hhhj��  hj��  ubj��  ]�(j7�  hs)��}�(hvKhwKhj��  hxh|j  K+hj��  hrj9  )��}�(hK	hK hj69  )��}�(hKhKhKhhhhh�h�hKh�hhhKh�hKh�Spear�h�ubhKh�h �j�  �h!K h"�hj��  h-KhKh.K hK hfj>9  )��}�(h�h�hKhhhKh.K
h�hhhj�  hhmubj�  G?�������h\KhDNj�  Nhd]�hFKdhHKh�Goblin Lancer�hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  KhqjE�  j�  j<9  )��}�(h�h�hKhhhKh.Kh�hhhj��  hj��  ubj��  ]�(j7�  jE�  hs)��}�(hvKhwK
hj��  hxh|j  K#hj��  hrj9  )��}�(hKhK hj29  )��}�(hKhKhKhhhhh�h�hKh�hhhKh�hKhj(�  h�ubhKh�h �j�  �h!K h"�hj��  h-KhKh.K hK hfj>9  )��}�(h�h�hKhhhKh.K
h�hhhj�  hhmubj�  G        h\KhDNj�  Nhd]�hFKdhHKhj,�  hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  KhqjU�  j�  j<9  )��}�(h�h�hKhhhKh.Kh�hhhj��  hj��  ubj��  ]�(j7�  jU�  ej�  Nj�  �hKububhs)��}�(hvKhwKhjρ  hxh|j  K.hj��  hrj�8  )��}�(hKhK hh�Mace���)��}�(hKhKhKhhhj�  h�h�hKh�hhhKh�hKh�Mace�h�ubhKh�h �j�  �h!K h"�hjρ  h-K	hKh.K hK hfjB9  )��}�(h�h�hKhhhKh.Kh�hhhj�  hhmubj�  G        h\KhDNj�  Nhd]�hFKdhHKh�Goblin Stonewall�hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqjc�  j�  j@9  )��}�(h�h�hKhhhK7h.K2h�hhh�Iron Breastplate�hj��  ubj��  ]�(jE�  jc�  ej�  j*9  )��}�(hKhKhhhj�  h�h�h�h�hhhKh.Kh�hK h�Iron Shield�hK ubj�  �hKububej�  j,9  )��}�(hKhKhhh�0H�h�h�h�h�hhhKh.Kh�hK h�Buckler�hK ubj�  �hKububjU�  jc�  ej�  Nj�  �hKububKjE�  Khs)��}�(hvKhwKhj́  hxh|j  K+h�Chest�hr�Features.Features��Chest���)��}�(hqj}�  hO]�(jD9  )��}�(h�h�hKhhhK#h.K#h�hhh�Chain Shirt�hj��  ubj89  )��}�(hKhKhKhhhj�  h�h�hKh�hhhKh�hKh�Dagger�h�ubj.9  )��}�(hKhKhhhj�  h�h�h�h�hhhKh.Kh�hK hj�  hK ubhQ�
Gold_Coins���)��}�(h��coins�Kh�h�$�h]�(K�K�Keh�
Gold Coins�hhYubehj́  h]�(KQKOKehj�  ububK	hs)��}�(hvKhwK	hhhxh|j  K(hjڂ  hrj.9  )��}�(hqj��  hKhKhhhj�  h�h�h�h�hhhKh.Kh�hK hj�  hK ububK
jU�  Kjc�  Khs)��}�(hvK"hwKhjӁ  hxh|j  KAh�	Stairs Up�hr�Features.Stairs��StairUp���)��}�(hqj��  hvK"hwJ����hxh|j  KA�moveCost�Kh�Stairs�hrNububKhtKhs)��}�(hvK5hwKhhWhxh|j  K=hj4�  hrhS)��}�(hVKh�h�hhWhqj��  hhhhXhhYububKhs)��}�(hvK7hwKhjρ  hxh|j  K=hj��  hrj�8  )��}�(hKhK hjh�  )��}�(hKhKhKhhhj�  h�h�hKh�hhhKh�hKhjk�  h�ubhKh�h �j�  �h!K h"�hjρ  h-KhKh.K hK hfjB9  )��}�(h�h�hKhhhKh.Kh�hhhj�  hhmubj�  G        h\KhDNj�  Nhd]�hFKdhHKhjo�  hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqj��  j�  j@9  )��}�(h�h�hKhhhK7h.K2h�hhhjt�  hj��  ubj��  ]�j�  j*9  )��}�(hKhKhhhj�  h�h�h�h�hhhKh.Kh�hK hjx�  hK ubj�  �hKububKhs)��}�(hvK7hwKhj��  hxh|j  K@hj��  hrj9  )��}�(hKhK hj29  )��}�(hKhKhKhhhhh�h�hKh�hhhKh�hKhj(�  h�ubhKh�h �j�  �h!K h"�hj��  h-KhKh.K hK hfj>9  )��}�(h�h�hKhhhKh.K
h�hhhj�  hhmubj�  G        h\KhDNj�  Nhd]�hFKdhHKhj,�  hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqj��  j�  j<9  )��}�(h�h�hKhhhKh.Kh�hhhj��  hj��  ubj��  ]�j�  Nj�  �hKububKhs)��}�(hvK;hwKhj́  hxh|j  Khj�  hrj��  )��}�(hqjǃ  hO]�(j*9  )��}�(hKhKhhhj�  h�h�h�h�hhhKh.Kh�hK hjx�  hK ubj*9  )��}�(hKhKhhhj�  h�h�h�h�hhhKh.Kh�hK hjx�  hK ubhi)��}�(h�h�hKhhhKh.Kh�hhhhlhhmubj��  )��}�(h�j��  Kh�hj��  hj��  hj��  hhYubehj́  hj��  hj�  ububKhs)��}�(hvK<hwKhj��  hxh|j  Khj��  hrj9  )��}�(hKhK hj29  )��}�(hKhKhKhhhhh�h�hKh�hhhKh�hKhj(�  h�ubhKh�h �j�  �h!K h"�hj��  h-KhKh.K hK hfj>9  )��}�(h�h�hKhhhKh.K
h�hhhj�  hhmubj�  G        h\KhDNj�  Nhd]�hFKdhHKhj,�  hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqjԃ  j�  j<9  )��}�(h�h�hKhhhKh.Kh�hhhj��  hj��  ubj��  ]�j�  Nj�  �hKububKhs)��}�(hvK=hwKhj��  hxh|j  Khj��  hrj"9  )��}�(hK	hK hj09  )��}�(hKhKhKhhhj�  h�h�hKh�hhhKh�hKhj�  h�ubhKh�h �j�  �h!K h"�hj��  h-KhKh.K hK hfj>9  )��}�(h�h�hKhhhKh.K
h�hhhj�  hhmubj�  G?��Q�h\KhDNj�  Nhd]�hFKdhHKhj�  hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqj�  j�  j<9  )��}�(h�h�hKhhhKh.Kh�hhhj��  hj��  ubj��  ]�j�  Nj�  �hKububKhs)��}�(hvK=hwKhj��  hxh|j  Khj��  hrj9  )��}�(hK
hK hj49  )��}�(hKhKhKhhhhh�h�hKh�hhhKh�hKhj݂  h�ubhKh�h �j�  �h!Kh"�hj��  h-KhKh.K hK hfhi)��}�(h�h�hKhhhKh.Kh�hhhhlhhmubj�  G?�      h\KhDNj�  Nhd]�hFKdhHKhj�  hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqj��  j�  j<9  )��}�(h�h�hKhhhKh.Kh�hhhj��  hj��  ubj��  ]�j�  Nj�  �hKububKhs)��}�(hvK=hwKhhWhxh|j  Khj4�  hrhS)��}�(hVKh�h�hhWhqj��  hhhhXhhYububKhs)��}�(hvK>hwKhj��  hxh|j  Khj��  hrj9  )��}�(hK
hK hj49  )��}�(hKhKhKhhhhh�h�hKh�hhhKh�hKhj݂  h�ubhKh�h �j�  �h!Kh"�hj��  h-KhKh.K hK hfhi)��}�(h�h�hKhhhKh.Kh�hhhhlhhmubj�  G?�      h\KhDNj�  Nhd]�hFKdhHKhj�  hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqj�  j�  j<9  )��}�(h�h�hKhhhKh.Kh�hhhj��  hj��  ubj��  ]�j�  Nj�  �hKububKhs)��}�(hvK>hwKhjρ  hxh|j  Khj��  hrj�8  )��}�(hKhK hjh�  )��}�(hKhKhKhhhj�  h�h�hKh�hhhKh�hKhjk�  h�ubhKh�h �j�  �h!K h"�hjρ  h-KhKh.K hK hfjB9  )��}�(h�h�hKhhhKh.Kh�hhhj�  hhmubj�  G        h\KhDNj�  Nhd]�hFKdhHKhjo�  hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqj�  j�  j@9  )��}�(h�h�hKhhhK7h.K2h�hhhjt�  hj��  ubj��  ]�j�  j*9  )��}�(hKhKhhhj�  h�h�h�h�hhhKh.Kh�hK hjx�  hK ubj�  �hKububKhs)��}�(hvK?hwKhhhxh|j  Khjڂ  hrj,9  )��}�(hqj �  hKhKhhhj{�  h�h�h�h�hhhKh.Kh�hK hj|�  hK ububKhs)��}�(hvK?hwKhhWhxh|j  K'hj4�  hrhS)��}�(hVKh�h�hhWhqj$�  hhhhXhhYububKhs)��}�(hvK@hwKhjρ  hxh|j  K$hj��  hrj�8  )��}�(hKhK hjh�  )��}�(hKhKhKhhhj�  h�h�hKh�hhhKh�hKhjk�  h�ubhKh�h �j�  �h!K h"�hjρ  h-K	hKh.K hK hfjB9  )��}�(h�h�hKhhhKh.Kh�hhhj�  hhmubj�  G        h\KhDNj�  Nhd]�hFKdhHKhjo�  hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqj(�  j�  j@9  )��}�(h�h�hKhhhK7h.K2h�hhhjt�  hj��  ubj��  ]�j�  j*9  )��}�(hKhKhhhj�  h�h�h�h�hhhKh.Kh�hK hjx�  hK ubj�  �hKububKhs)��}�(hvK@hwKhj��  hxh|j  K%hj��  hrj9  )��}�(hKhK hj29  )��}�(hKhKhKhhhhh�h�hKh�hhhKh�hKhj(�  h�ubhKh�h �j�  �h!K h"�hj��  h-KhKh.K hK hfj>9  )��}�(h�h�hKhhhKh.K
h�hhhj�  hhmubj�  G        h\KhDNj�  Nhd]�hFKdhHKhj,�  hJK hO]�hCK h]]�hj�  j�  Nh`K j��  K(j�  K j�  NhE�hcNhnKho�j�  Khqj8�  j�  j<9  )��}�(h�h�hKhhhKh.Kh�hhhj��  hj��  ubj��  ]�j�  Nj�  �hKububKhs)��}�(hvKAhwKhj�  hxh|j  K"h�Stairs Down�hrj��  �	StairDown���)��}�(hqjF�  hrNhwJ����hxh|hvKAj��  Khj��  j  K"ububu�consumeList�]�(hSjЂ  j҂  jԂ  jւ  eh�
1B: Forest��djikstra_Player_Adj�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K%K$K#K"K!Ne]�(NK_K^K]K\NNKYKXKWKVKUKTKSKRKQKPKOKNKMNKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$K#K$K#NK!K Ne]�(NK^K]K\K[KZNKXKWKVKUKTNNKQNKOKNKMKLKKKJNKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K#K"K!K KNe]�(NK]K\K[NKYKXKWKVNKTKSKRKQKPNKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K"K!K KKNe]�(NK\K[KZNKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,NK*K)NK'K&K%K$K#K"K!K NK KKKNe]�(NK[KZKYKXKWKVKUKTKSKRKQKPKONKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(K'NK%K$K#K"K!K KK KNKKNe]�(NKZKYKXKWKVKUKTKSKRKQNKOKNKMKLKKKJNKHNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*NK(K'K&K%K$K#K"K!K KKKKKKKNe]�(NKYKXNKVKUKTKSKRKQKPKOKNNKLKKNKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&NK$K#NK!K KKKKKKKKNe]�(NKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKGNKCKBNNK?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"NK KKKKKNKKKNe]�(NKWKVKUKTKSKTKSNKOKNKMKLKKNKIKHKGKFKENKCNKAK@K?K>K=K<NK:K9K8K7K6K5K4K3K2K1K0K/K.NK,K+K*K)K(K'K&K%K$K#K"K!K KKKNKKKKKKNe]�(NKVKUNKSKRKSNKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?NK=K<K;K:K9K8NNK5K4K3K2K1K0K/K.K-K,NK*K)K(K'K&K%K$K#K"K!K KKKNKKKKKKKNe]�(NKUKTKSKRKQNKOKNKMKLKKKLNKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKNKKKKNe]�(NKTKSKRKQKPKOKNKMNKKKJNKHNKFKEKDKCKBKAK@K?NK=K<K;K:K9K8K7K6K5NK3K2K1K0K/K.K-K,K+K*K)K(K'NNK$K#K"K!K KKKKKKKKKKKKKNe]�(NKSKRKQKPKOKNKMKLKKKJKINKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K KKKKKKKKKKKKKKNe]�(NKRKQKPKOKNKMKLKKKJKIKHKGKFNKDKCKBKAK@NK>K=K<K;K:K9K8K7NNK4K3NK1K0K/K.K-K,K+K*K)K(K'K&K%K$NK"K!K KKKKKKNKKKKKKKKNe]�(NKQKPKOKNKMNKMNKIKHKGKFKEKDKCKBKAK@K?K>NK<K;K:NK8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K KKKKKKKNKKKKKKKKNe]�(NKPKONKMKLKKKLKKKJKINKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!NKKKKKKKKKNKKKKKKKNe]�(NKOKNKMKLKKKJKKKLKKKJNKDKCKBKAKBNK>K=K<K;K:NK8NK6NK4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKNe]�(NKNKMKLKKKJKIKJKKNNKDNKBKAK@NK>K=K<K;K:K9NK7K6K5K4NK2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKNe]�(NKMKLKKKJKIKHNNKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5NK3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKNe]�(NKLKKKJNKHKGKFKEKDNKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKNe]�(NKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/NK-K,NK*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKNe]�(NKLKKKJKINKGKFNKDKCKBKAK@K?K>K=K<K;K:NK6K5K4K3K2NK0K/K.NK,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKNe]�(NKMNKKKJKINKGKFKEKDNKBKAK@K?K>K=K<K;NK5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKK
Ne]�(NKLKKKJKIKHKGKFKEKDNKBKAK@K?K>K=K<K;K:NK6K5K4K3NK1K0NK,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKK
K	Ne]�(NKKKJKIKHKGKFKEKDKCKBNK@NNK=K<K;K:K9K8K7K6NK2K1K0K/K.K-K,K+K*K)NNNNNNNNNNNNNNNNKKKKKKKKNKKKNKK
K	KNe]�(NKJKIKHKGKFNKDKCKBKAK@K?K>K=K<K;NK9K8K7K6K5NK3K2K1K0K/K.K-K,K+K*NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NKKKKKKKKKNKK
K	K
K	KKNe]�(NKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4NK2K1K0K/K.K-K,K+K*K)NK+K,K-K.K/K0K1K2K3K4K5K6K7K8NKKKKKKKKKKK
K	KK	KKKNe]�(NKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NK8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7NKKKKKKKKKK
K	KKKKKKNe]�(NKIKHKGKFKENNNKAK@K?NK=NK;K:NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK+K,K-K.K/K0K1K2K3K4K5K6K7K8NKKKKKKKKNK	KKKKKKKNe]�(NKHKGKFKEKDKCNKAK@K?K>K=K<K;K:K9K8K7NK3K2K1K0K/K.K-K,K+K*K)K(K'K&NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NKKKKKKKK
K	KKKKKKKKNe]�(NKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2NK.K-K,K+K*K)K(K'K&K%NK-K.K/K0K1K2K3K4K5K6K7K8K9K:NKKKKKKK
K	KKKKKKNKKNe]�(NKFNKDKCNKAK@K?NK=K<K;K:K9K8K7K6K5K4K3K2K1K0NK,K+K*K)K(K'K&K%K$NNNNNNNNNNNNNNNNKKKKKKKK
NKKKKNKK KNe]�(NKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK$K#K"K!K KKKKKKKKKKKKKKNNKKKKKNKKKKKK KK Ne]�(NKFNKDNKBKAK@K?K>NK<K;K:K9K8NK4K3K2K1K0K/K.K-K,NK*NK(NK&K%K$K#K"K!K KKKKKKKKKKKKKKKKKNKKNKKKKKKK KNe]�(NKGKFKEKDKCNKAK@K?NK;K:K9K8K7K6K5K4K3K2NK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKNKKKKKNKKNe]�(NKHNNKCKBNK@K?K>K=K<NK8K7K6K5K4K3K2K1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKNKK
K	KKKKKKKKNe]�(NKGKFKENKAK@K?K>K=K<K;K:K9K8K7K6K5NNK2NK0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K KKKKKKKKKKKNKKKKKKKNK	KNNKKKKNe]�(NKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4NNK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKNKK
K	KKKKKKNe]�(NKGKFKEKDKCKBKAK@K?NK=K<K;K:K9K8NK4K3K2K1K0NK.K-K,K+K*K)NK'K&K%K$K#K"K!K KKKKKKKKKKKKNKKKKKKKKK
K	KKKKKNe]�(NKHKGKFKEKDNKBKAK@K?K>NK:K9K8K7K6K5K4K3K2K1K0K/K.K-NK+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKNKKKKKKKKKNK	KKKKNe]�(NKIKHNKDKCKBKAK@K?K>K=K<K;NK9K8NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"NK NKKKKKKKKKKKKKKKKKKKKK
K	KKKNe]�(NKHKGKFKEKDKCNKANK?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#NK!K KKKKNKKNKKKKKKKKKKKKKK
K	KK	Ne]�(NKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK8K7K6K5K4K3NK1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!NKKKKKKKKKNKKKKNKKKKKKK
K	K
Ne]�(NKJKIKHKGKFKEKDKCKBKAK@K?K>K=NK;K:K9NK7K6K5NK3K2K1K0K1NK-K,K+K*K)NNK&NK$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
KNe]�(NKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK8K7K6NK4K3K2K1K0K/K.NK,K+K*K)K(K'K(NK$K#K"K!K KKKNKKKKKNKKNKKKKKKKKKNe]�(NKLKKKJKIKHKGKFKENKCKBKAK@NNNNK;K:K9K8K7K6K5NK3K2K1K0K/K.K-K,K+K*K)K(K)NK%K$K#K"K!K KKKKKNKKKKKKKKKKKKKKKNe]�(NKMKLKKKJKIKHNKFNKDKCKBKAK@K?K>K=K<K;K:NK8K7K6K7NK3K2K1NK/K.K-K,K+K*K)K(K'K&K%K$K#K"NK KKNKKNKKKNKKKKKKKKKKNe]�(NKNKMKLKKNKINKGKFKEKDKCKBKAK@K?K>K=NK;K:K9K8K7K6K5K4K3K2NK0K/K.K-K,K+K*K)K(K'K&K%NK#K"K!K KKKKKKKKNKKKKKKKKKKNe]�(NKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5NK3K2K1NK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKNe]�(NKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%NK#K"K!K KKKKKKKKKKKKKKKKKNe]�(NKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKNe]�(NKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKNe]�(NKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)NK'K&K%K$K#K"K!K KKKKKKKKKKKKKKNe]�(NKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;NK9K8NK6K5K4K3K2K1K0K/K.K-K,K+K*NK(K'NK%K$K#K"K!K KKKKKKKKKKKKKNe]�(NKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,NK*K)K(NK&K%K$K#K"K!K KKKKKKKKKKKKNe]�(NKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*NK(K'K&K%K$K#K"K!K KKKKKKKKKKKNe]�(NKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7NNNNNNNNK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKNe]�(NKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8NK>K?K@KAKBKCNK/K.K-K,K+K*K)K(NK&K%NK#K"K!K KKKKKKKKKNe]�(NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK=K>K?K@KAKBNK0K/K.K-K,K+K*K)K(K'K&NK$K#K"K!K KKKKKKKKNe]�(NKZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K;K<K=K>K?K@KANK1K0K/K.K-K,K+K*K)K(K'K(NK$K#NK!K KKKKKKKNe]�(NK[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;NK=K>K?K@KAKBNK2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K!K KKKKKKNe]�(NK\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NK>K?K@KAKBKCNK3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K KKKKKNe]�(NK]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=NK?K@KAKBKCKDNK4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K!K KKKKNe]�(NK^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K?NNNNNNNK5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKNe]�(NK_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KK Ne]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�cLevel�Kubj  KAh�Player�hrhubj�  j:9  )��}�(h�h�hKhhhKh.Kh�hhh�Cloth Shirt�hj��  ubj�  h�Tome���)��}�(hK hKhKhhhj{�  h�h�hKh�hhhKh�hK h�Tome�h�ubj�  �j�  Nub.