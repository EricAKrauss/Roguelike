��      �__main__��Game���)��}�(�width�K#�loadRequest���yConst�KK�turn�K�	thePlayer��Player�h
��)��}�(�	sightDist�K�accuracy�K �	rightHand��Items.Weapons��Staff���)��}�(�armorPen�K�level�K�range�K�color�]�(K�K�K�e�type��2H��
equippable���addPower���magPower�K�
usesArrows���char��?��weight�K�	throwable���power�K�name��Staff��
consumable��ubhK�visible���canMove���arrows�K �invertColor��h!�@��skillLevels�}�(�6�K �2�K �3�K �7�K �1�K �5�K �4�K u�gold�K hK�armorVal�K hK �rightScroll�N�skillPoints�Kh%K�
baseHealth�K��skills�}�(h0�	Abilities��Flash_Freeze���h1h>�Shocking_Grasp���h2h>�Fireball���h3h>�Arcane_Reservoir���h4h>�Blink���h5h>�Wall_of_Force���h6h>�Lightning_Bolt���u�
healthTemp�K �	rightRing�N�playerControlled���expNext�Kd�healthCurve�G?�      �	healthMax�K�h&�Kyle��dodge�K �Class��Player_Classes��Mage����items�]�(�Items.Consumables��	GreenHerb���)��}�(�healNum�Kh�h(�h!�+�hhh&�
Green Herb�h�
consumable�ubh])��}�(h`Kh�h(�h!hahhh&hbhhcube�
initiative�K�effects�]�h]�(KKYK�e�exp�K �
leftScroll�N�recalcTimer�K �leftRing�N�
hitEffects�]��helmet��Items.Armors��	Cloth_Hat���)��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&�	Cloth Hat�h�helmet�ub�health�K��
countering���	recalcMax�K �pObject��Object�h|��)��}�(�row�K"�ID�Kh!h-�pLevel��LevelTypes.LevelTypes��Wild���)��}�(�	decorList�]�(�LevelTypes.Decorations��Table���h��Firepit���h��Weapon_Rack���eh	h�master_Changed_Tiles�]�(]�(K!K@e]�(K K?e]�(KK>e]�(KK=e]�(KK<e]�(KK;e]�(KK:e]�(KK9e]�(K!KBe]�(K KCe]�(K!K@e]�(K K?e]�(KK>e]�(KK=e]�(KK<e]�(KK;e]�(KK:e]�(KK9e]�(K!KBe]�(K KCe]�(K!K@e]�(K K?e]�(KK>e]�(KK=e]�(KK<e]�(KK;e]�(KK:e]�(KK9e]�(K!KBe]�(K KCe]�(K!K@e]�(K K?e]�(K K>e]�(KK=e]�(KK<e]�(KK;e]�(KK:e]�(KK9e]�(K!KBe]�(K!KCe]�(K!K@e]�(K!K?e]�(K!KBe]�(K!KCe]�(K!K@e]�(K!K?e]�(K!KBe]�(K!KCe]�(K!K@e]�(K!K?e]�(K"KBe]�(K!KCe]�(K"K@e]�(K!K?e]�(K"KBe]�(K!KCe]�(K"K@e]�(K!K?e]�(K"KBe]�(K!KCe]�(K"K@e]�(K!K?e]�(K"KBe]�(K"KCe]�(K"K@e]�(K"K?e]�(K!K>e]�(K!K=e]�(K!K<e]�(K!K;e]�(K!K:e]�(K"KBe]�(K"KCe]�(K"K@e]�(K"K?e]�(K"K>e]�(K"K=e]�(K"K<e]�(K!K;e]�(K!K:e]�(K"KBe]�(K"KCe]�(K"K@e]�(K"K?e]�(K"K>e]�(K"K=e]�(K"K<e]�(K"K;e]�(K"K:e]�(K"KBe]�(K"KCe]�(K"K@e]�(K"K?e]�(K"K>e]�(K"K=e]�(K"K<e]�(K#K;e]�(K#K:e]�(K"KBe]�(K"KCe]�(K"K@e]�(K"K?e]�(K#K>e]�(K#K=e]�(K#K<e]�(K#K;e]�(K#K:e]�(K"KBe]�(K"KCe]�(K"K@e]�(K#K?e]�(K#K>e]�(K#K=e]�(K#K<e]�(K$K;e]�(K$K:e]�(K"KBe]�(K"KCe]�(K"K@e]�(K#K?e]�(K#K>e]�(K#K=e]�(K$K<e]�(K$K;e]�(K$K:e]�(K"KBe]�(K#KCe]�(K"K@e]�(K#K?e]�(K#K>e]�(K$K=e]�(K$K<e]�(K%K;e]�(K%K:e]�(K%K9e]�(K"KBe]�(K#KCe]�(K#K@e]�(K#K?e]�(K$K>e]�(K$K=e]�(K%K<e]�(K%K;e]�(K&K:e]�(K"KBe]�(K#KCe]�(K#K@e]�(K#K?e]�(K$K>e]�(K$K=e]�(K%K<e]�(K&K;e]�(K&K:e]�(K#KBe]�(K#KCe]�(K#K@e]�(K#K?e]�(K$K>e]�(K%K=e]�(K%K<e]�(K&K;e]�(K'K:e]�(K'K9e]�(K#KBe]�(K#KCe]�(K#K@e]�(K$K?e]�(K$K>e]�(K%K=e]�(K&K<e]�(K'K;e]�(K'K:e]�(K(K9e]�(K#KBe]�(K#KCe]�(K#K@e]�(K$K?e]�(K%K>e]�(K%K=e]�(K&K<e]�(K'K;e]�(K(K:e]�(K)K9e]�(K#KBe]�(K$KCe]�(K#K@e]�(K$K?e]�(K%K>e]�(K&K=e]�(K#KBe]�(K$KCe]�(K#K@e]�(K$K?e]�(K%K>e]�(K&K=e]�(K#KBe]�(K$KCe]�(K!K@e]�(K K?e]�(KK>e]�(KK=e]�(KK<e]�(KK;e]�(KK:e]�(KK9e]�(K#K@e]�(K$K?e]�(K%K>e]�(K&K=e]�(K!K@e]�(K K?e]�(KK>e]�(KK=e]�(KK<e]�(KK;e]�(KK;e]�(K#K@e]�(K$K?e]�(K%K>e]�(K&K=e]�(K!K@e]�(K K?e]�(KK>e]�(KK>e]�(KK=e]�(KK<e]�(KK;e]�(K#K@e]�(K$K?e]�(K%K?e]�(K&K>e]�(K!K@e]�(K K?e]�(KK?e]�(KK>e]�(KK=e]�(KK<e]�(KK<e]�(KK;e]�(K#K@e]�(K$K@e]�(K!K@e]�(K K@e]�(K#K@e]�(K$K@e]�(K!K@e]�(K K@e]�(K#K@e]�(K$K@e]�(K!K@e]�(K K@e]�(K#KAe]�(K$K@e]�(K!KAe]�(K#KAe]�(K$K@e]�(K!KAe]�(K#KAe]�(K$K@e]�(K!KAe]�(K#KAe]�(K$KAe]�(K%K@e]�(K&K@e]�(K'K@e]�(K(K@e]�(K)K?e]�(K*K?e]�(K!KAe]�(K#KAe]�(K$KAe]�(K%KAe]�(K&K@e]�(K'K@e]�(K(K@e]�(K)K@e]�(K*K@e]�(K!KAe]�(K#KAe]�(K$KAe]�(K%KAe]�(K&KAe]�(K'KAe]�(K(KAe]�(K)K@e]�(K*K@e]�(K!KAe]�(K#KAe]�(K$KAe]�(K%KAe]�(K&KAe]�(K'KAe]�(K(KAe]�(K)KAe]�(K*KAe]�(K!KAe]�(K#KAe]�(K$KAe]�(K%KAe]�(K&KAe]�(K'KAe]�(K(KAe]�(K)KBe]�(K*KBe]�(K!KAe]�(K#KAe]�(K$KAe]�(K%KAe]�(K&KBe]�(K'KBe]�(K(KBe]�(K)KBe]�(K*KBe]�(K!KAe]�(K#KAe]�(K$KAe]�(K%KBe]�(K&KBe]�(K'KBe]�(K(KBe]�(K)KCe]�(K!KAe]�(K#KAe]�(K$KBe]�(K%KBe]�(K&KBe]�(K'KCe]�(K!KAe]�(K#KAe]�(K$KBe]�(K%KBe]�(K&KCe]�(K!KBe]�(K KBe]�(KKCe]�(K#KAe]�(K$KBe]�(K%KBe]�(K&KCe]�(K!KBe]�(K KBe]�(KKCe]�(K#KBe]�(K$KBe]�(K%KCe]�(K!KBe]�(K KBe]�(KKCe]�(K#KBe]�(K$KBe]�(K%KCe]�(K!KBe]�(K KCe]�(K#KBe]�(K$KBe]�(K%KCe]�(K!KBe]�(K KCe]�(K#KBe]�(K$KCe]�(K!KBe]�(K KCe]�(K#KBe]�(K$KCe]�(K!KBe]�(K KCe]�(K#KBe]�(K$KCee�
stairsDown�]�(KAK"e�Tiles�}�(K }�(K �Tile�j  ��)��}�(h�K �Objects�]�h�h��col�K ubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubK	j	  )��}�(h�K j  ]�h�h�j  K	ubK
j	  )��}�(h�K j  ]�h�h�j  K
ubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubK j	  )��}�(h�K j  ]�h�h�j  K ubK!j	  )��}�(h�K j  ]�h�h�j  K!ubK"j	  )��}�(h�K j  ]�h�h�j  K"ubK#j	  )��}�(h�K j  ]�h�h�j  K#ubK$j	  )��}�(h�K j  ]�h�h�j  K$ubK%j	  )��}�(h�K j  ]�h�h�j  K%ubK&j	  )��}�(h�K j  ]�h�h�j  K&ubK'j	  )��}�(h�K j  ]�h�h�j  K'ubK(j	  )��}�(h�K j  ]�h�h�j  K(ubK)j	  )��}�(h�K j  ]�h�h�j  K)ubK*j	  )��}�(h�K j  ]�h�h�j  K*ubK+j	  )��}�(h�K j  ]�h�h�j  K+ubK,j	  )��}�(h�K j  ]�h�h�j  K,ubK-j	  )��}�(h�K j  ]�h�h�j  K-ubK.j	  )��}�(h�K j  ]�h�h�j  K.ubK/j	  )��}�(h�K j  ]�h�h�j  K/ubK0j	  )��}�(h�K j  ]�h�h�j  K0ubK1j	  )��}�(h�K j  ]�h�h�j  K1ubK2j	  )��}�(h�K j  ]�h�h�j  K2ubK3j	  )��}�(h�K j  ]�h�h�j  K3ubK4j	  )��}�(h�K j  ]�h�h�j  K4ubK5j	  )��}�(h�K j  ]�h�h�j  K5ubK6j	  )��}�(h�K j  ]�h�h�j  K6ubK7j	  )��}�(h�K j  ]�h�h�j  K7ubK8j	  )��}�(h�K j  ]�h�h�j  K8ubK9j	  )��}�(h�K j  ]�h�h�j  K9ubK:j	  )��}�(h�K j  ]�h�h�j  K:ubK;j	  )��}�(h�K j  ]�h�h�j  K;ubK<j	  )��}�(h�K j  ]�h�h�j  K<ubK=j	  )��}�(h�K j  ]�h�h�j  K=ubK>j	  )��}�(h�K j  ]�h�h�j  K>ubK?j	  )��}�(h�K j  ]�h�h�j  K?ubK@j	  )��}�(h�K j  ]�h�h�j  K@ubKAj	  )��}�(h�K j  ]�h�h�j  KAubKBj	  )��}�(h�K j  ]�h�h�j  KBubKCj	  )��}�(h�K j  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�K ah�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�Kah�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�Kah�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK	}�(K j	  )��}�(h�K	j  ]�h�h�j  K ubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubK	j	  )��}�(h�K	j  ]�h�h�j  K	ubK
j	  )��}�(h�K	j  ]�h�h�j  K
ubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubKj	  )��}�(h�K	j  ]�h�h�j  KubK j	  )��}�(h�K	j  ]�h�h�j  K ubK!j	  )��}�(h�K	j  ]�h�h�j  K!ubK"j	  )��}�(h�K	j  ]�h�h�j  K"ubK#j	  )��}�(h�K	j  ]�h�h�j  K#ubK$j	  )��}�(h�K	j  ]�h�h�j  K$ubK%j	  )��}�(h�K	j  ]�h�h�j  K%ubK&j	  )��}�(h�K	j  ]�h�h�j  K&ubK'j	  )��}�(h�K	j  ]�h�h�j  K'ubK(j	  )��}�(h�K	j  ]�h�h�j  K(ubK)j	  )��}�(h�K	j  ]�h�h�j  K)ubK*j	  )��}�(h�K	j  ]�h�h�j  K*ubK+j	  )��}�(h�K	j  ]�h�h�j  K+ubK,j	  )��}�(h�K	j  ]�h�h�j  K,ubK-j	  )��}�(h�K	j  ]�h�h�j  K-ubK.j	  )��}�(h�K	j  ]�h�h�j  K.ubK/j	  )��}�(h�K	j  ]�h�h�j  K/ubK0j	  )��}�(h�K	j  ]�h�h�j  K0ubK1j	  )��}�(h�K	j  ]�h�h�j  K1ubK2j	  )��}�(h�K	j  ]�h�h�j  K2ubK3j	  )��}�(h�K	j  ]�h�h�j  K3ubK4j	  )��}�(h�K	j  ]�h�h�j  K4ubK5j	  )��}�(h�K	j  ]�h�h�j  K5ubK6j	  )��}�(h�K	j  ]�h�h�j  K6ubK7j	  )��}�(h�K	j  ]�h�h�j  K7ubK8j	  )��}�(h�K	j  ]�h�h�j  K8ubK9j	  )��}�(h�K	j  ]�h�h�j  K9ubK:j	  )��}�(h�K	j  ]�h�h�j  K:ubK;j	  )��}�(h�K	j  ]�h�h�j  K;ubK<j	  )��}�(h�K	j  ]�h�h�j  K<ubK=j	  )��}�(h�K	j  ]�h�h�j  K=ubK>j	  )��}�(h�K	j  ]�h�h�j  K>ubK?j	  )��}�(h�K	j  ]�h�h�j  K?ubK@j	  )��}�(h�K	j  ]�h�h�j  K@ubKAj	  )��}�(h�K	j  ]�h�h�j  KAubKBj	  )��}�(h�K	j  ]�h�h�j  KBubKCj	  )��}�(h�K	j  ]�h�h�j  KCubuK
}�(K j	  )��}�(h�K
j  ]�h�h�j  K ubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubK	j	  )��}�(h�K
j  ]�h�h�j  K	ubK
j	  )��}�(h�K
j  ]�h�h�j  K
ubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubKj	  )��}�(h�K
j  ]�h�h�j  KubK j	  )��}�(h�K
j  ]�h�h�j  K ubK!j	  )��}�(h�K
j  ]�h�h�j  K!ubK"j	  )��}�(h�K
j  ]�h�h�j  K"ubK#j	  )��}�(h�K
j  ]�h�h�j  K#ubK$j	  )��}�(h�K
j  ]�h�h�j  K$ubK%j	  )��}�(h�K
j  ]�h�h�j  K%ubK&j	  )��}�(h�K
j  ]�h�h�j  K&ubK'j	  )��}�(h�K
j  ]�h�h�j  K'ubK(j	  )��}�(h�K
j  ]�h�h�j  K(ubK)j	  )��}�(h�K
j  ]�h�h�j  K)ubK*j	  )��}�(h�K
j  ]�h�h�j  K*ubK+j	  )��}�(h�K
j  ]�h�h�j  K+ubK,j	  )��}�(h�K
j  ]�h�h�j  K,ubK-j	  )��}�(h�K
j  ]�h�h�j  K-ubK.j	  )��}�(h�K
j  ]�h�h�j  K.ubK/j	  )��}�(h�K
j  ]�h�h�j  K/ubK0j	  )��}�(h�K
j  ]�h�h�j  K0ubK1j	  )��}�(h�K
j  ]�h�h�j  K1ubK2j	  )��}�(h�K
j  ]�h�h�j  K2ubK3j	  )��}�(h�K
j  ]�h�h�j  K3ubK4j	  )��}�(h�K
j  ]�h�h�j  K4ubK5j	  )��}�(h�K
j  ]�h�h�j  K5ubK6j	  )��}�(h�K
j  ]�h�h�j  K6ubK7j	  )��}�(h�K
j  ]�h�h�j  K7ubK8j	  )��}�(h�K
j  ]�h�h�j  K8ubK9j	  )��}�(h�K
j  ]�h�h�j  K9ubK:j	  )��}�(h�K
j  ]�h�h�j  K:ubK;j	  )��}�(h�K
j  ]�h�h�j  K;ubK<j	  )��}�(h�K
j  ]�h�h�j  K<ubK=j	  )��}�(h�K
j  ]�h�h�j  K=ubK>j	  )��}�(h�K
j  ]�h�h�j  K>ubK?j	  )��}�(h�K
j  ]�h�h�j  K?ubK@j	  )��}�(h�K
j  ]�h�h�j  K@ubKAj	  )��}�(h�K
j  ]�h�h�j  KAubKBj	  )��}�(h�K
j  ]�h�h�j  KBubKCj	  )��}�(h�K
j  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�Kah�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�Kah�h�j  K5ubK6j	  )��}�(h�Kj  ]�Kah�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  �       KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�Kah�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�Kah�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�Kah�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�h�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�K	ah�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�h�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�h�j  K ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK	j	  )��}�(h�Kj  ]�h�h�j  K	ubK
j	  )��}�(h�Kj  ]�h�h�j  K
ubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubKj	  )��}�(h�Kj  ]�h�h�j  KubK j	  )��}�(h�Kj  ]�h�h�j  K ubK!j	  )��}�(h�Kj  ]�h�h�j  K!ubK"j	  )��}�(h�Kj  ]�h�h�j  K"ubK#j	  )��}�(h�Kj  ]�K
ah�h�j  K#ubK$j	  )��}�(h�Kj  ]�h�h�j  K$ubK%j	  )��}�(h�Kj  ]�h�h�j  K%ubK&j	  )��}�(h�Kj  ]�h�h�j  K&ubK'j	  )��}�(h�Kj  ]�h�h�j  K'ubK(j	  )��}�(h�Kj  ]�h�h�j  K(ubK)j	  )��}�(h�Kj  ]�h�h�j  K)ubK*j	  )��}�(h�Kj  ]�h�h�j  K*ubK+j	  )��}�(h�Kj  ]�h�h�j  K+ubK,j	  )��}�(h�Kj  ]�h�h�j  K,ubK-j	  )��}�(h�Kj  ]�h�h�j  K-ubK.j	  )��}�(h�Kj  ]�Kah�h�j  K.ubK/j	  )��}�(h�Kj  ]�h�h�j  K/ubK0j	  )��}�(h�Kj  ]�h�h�j  K0ubK1j	  )��}�(h�Kj  ]�h�h�j  K1ubK2j	  )��}�(h�Kj  ]�h�h�j  K2ubK3j	  )��}�(h�Kj  ]�h�h�j  K3ubK4j	  )��}�(h�Kj  ]�h�h�j  K4ubK5j	  )��}�(h�Kj  ]�h�h�j  K5ubK6j	  )��}�(h�Kj  ]�h�h�j  K6ubK7j	  )��}�(h�Kj  ]�h�h�j  K7ubK8j	  )��}�(h�Kj  ]�h�h�j  K8ubK9j	  )��}�(h�Kj  ]�h�h�j  K9ubK:j	  )��}�(h�Kj  ]�h�h�j  K:ubK;j	  )��}�(h�Kj  ]�h�h�j  K;ubK<j	  )��}�(h�Kj  ]�h�h�j  K<ubK=j	  )��}�(h�Kj  ]�h�h�j  K=ubK>j	  )��}�(h�Kj  ]�h�h�j  K>ubK?j	  )��}�(h�Kj  ]�h�h�j  K?ubK@j	  )��}�(h�Kj  ]�h�h�j  K@ubKAj	  )��}�(h�Kj  ]�h�h�j  KAubKBj	  )��}�(h�Kj  ]�h�h�j  KBubKCj	  )��}�(h�Kj  ]�h�h�j  KCubuK }�(K j	  )��}�(h�K j  ]�h�h�j  K ubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubK	j	  )��}�(h�K j  ]�h�h�j  K	ubK
j	  )��}�(h�K j  ]�h�h�j  K
ubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubKj	  )��}�(h�K j  ]�h�h�j  KubK j	  )��}�(h�K j  ]�h�h�j  K ubK!j	  )��}�(h�K j  ]�h�h�j  K!ubK"j	  )��}�(h�K j  ]�h�h�j  K"ubK#j	  )��}�(h�K j  ]�h�h�j  K#ubK$j	  )��}�(h�K j  ]�h�h�j  K$ubK%j	  )��}�(h�K j  ]�h�h�j  K%ubK&j	  )��}�(h�K j  ]�h�h�j  K&ubK'j	  )��}�(h�K j  ]�h�h�j  K'ubK(j	  )��}�(h�K j  ]�h�h�j  K(ubK)j	  )��}�(h�K j  ]�h�h�j  K)ubK*j	  )��}�(h�K j  ]�h�h�j  K*ubK+j	  )��}�(h�K j  ]�h�h�j  K+ubK,j	  )��}�(h�K j  ]�h�h�j  K,ubK-j	  )��}�(h�K j  ]�h�h�j  K-ubK.j	  )��}�(h�K j  ]�h�h�j  K.ubK/j	  )��}�(h�K j  ]�h�h�j  K/ubK0j	  )��}�(h�K j  ]�h�h�j  K0ubK1j	  )��}�(h�K j  ]�h�h�j  K1ubK2j	  )��}�(h�K j  ]�h�h�j  K2ubK3j	  )��}�(h�K j  ]�h�h�j  K3ubK4j	  )��}�(h�K j  ]�h�h�j  K4ubK5j	  )��}�(h�K j  ]�h�h�j  K5ubK6j	  )��}�(h�K j  ]�h�h�j  K6ubK7j	  )��}�(h�K j  ]�h�h�j  K7ubK8j	  )��}�(h�K j  ]�h�h�j  K8ubK9j	  )��}�(h�K j  ]�h�h�j  K9ubK:j	  )��}�(h�K j  ]�h�h�j  K:ubK;j	  )��}�(h�K j  ]�h�h�j  K;ubK<j	  )��}�(h�K j  ]�h�h�j  K<ubK=j	  )��}�(h�K j  ]�h�h�j  K=ubK>j	  )��}�(h�K j  ]�h�h�j  K>ubK?j	  )��}�(h�K j  ]�h�h�j  K?ubK@j	  )��}�(h�K j  ]�h�h�j  K@ubKAj	  )��}�(h�K j  ]�h�h�j  KAubKBj	  )��}�(h�K j  ]�h�h�j  KBubKCj	  )��}�(h�K j  ]�h�h�j  KCubuK!}�(K j	  )��}�(h�K!j  ]�h�h�j  K ubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubK	j	  )��}�(h�K!j  ]�h�h�j  K	ubK
j	  )��}�(h�K!j  ]�h�h�j  K
ubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubKj	  )��}�(h�K!j  ]�h�h�j  KubK j	  )��}�(h�K!j  ]�h�h�j  K ubK!j	  )��}�(h�K!j  ]�h�h�j  K!ubK"j	  )��}�(h�K!j  ]�h�h�j  K"ubK#j	  )��}�(h�K!j  ]�h�h�j  K#ubK$j	  )��}�(h�K!j  ]�h�h�j  K$ubK%j	  )��}�(h�K!j  ]�h�h�j  K%ubK&j	  )��}�(h�K!j  ]�h�h�j  K&ubK'j	  )��}�(h�K!j  ]�h�h�j  K'ubK(j	  )��}�(h�K!j  ]�h�h�j  K(ubK)j	  )��}�(h�K!j  ]�h�h�j  K)ubK*j	  )��}�(h�K!j  ]�h�h�j  K*ubK+j	  )��}�(h�K!j  ]�h�h�j  K+ubK,j	  )��}�(h�K!j  ]�h�h�j  K,ubK-j	  )��}�(h�K!j  ]�h�h�j  K-ubK.j	  )��}�(h�K!j  ]�h�h�j  K.ubK/j	  )��}�(h�K!j  ]�h�h�j  K/ubK0j	  )��}�(h�K!j  ]�h�h�j  K0ubK1j	  )��}�(h�K!j  ]�h�h�j  K1ubK2j	  )��}�(h�K!j  ]�h�h�j  K2ubK3j	  )��}�(h�K!j  ]�h�h�j  K3ubK4j	  )��}�(h�K!j  ]�h�h�j  K4ubK5j	  )��}�(h�K!j  ]�h�h�j  K5ubK6j	  )��}�(h�K!j  ]�h�h�j  K6ubK7j	  )��}�(h�K!j  ]�h�h�j  K7ubK8j	  )��}�(h�K!j  ]�h�h�j  K8ubK9j	  )��}�(h�K!j  ]�h�h�j  K9ubK:j	  )��}�(h�K!j  ]�h�h�j  K:ubK;j	  )��}�(h�K!j  ]�h�h�j  K;ubK<j	  )��}�(h�K!j  ]�h�h�j  K<ubK=j	  )��}�(h�K!j  ]�h�h�j  K=ubK>j	  )��}�(h�K!j  ]�h�h�j  K>ubK?j	  )��}�(h�K!j  ]�h�h�j  K?ubK@j	  )��}�(h�K!j  ]�h�h�j  K@ubKAj	  )��}�(h�K!j  ]�h�h�j  KAubKBj	  )��}�(h�K!j  ]�h�h�j  KBubKCj	  )��}�(h�K!j  ]�h�h�j  KCubuK"}�(K j	  )��}�(h�K"j  ]�h�h�j  K ubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubK	j	  )��}�(h�K"j  ]�h�h�j  K	ubK
j	  )��}�(h�K"j  ]�h�h�j  K
ubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubKj	  )��}�(h�K"j  ]�h�h�j  KubK j	  )��}�(h�K"j  ]�h�h�j  K ubK!j	  )��}�(h�K"j  ]�h�h�j  K!ubK"j	  )��}�(h�K"j  ]�h�h�j  K"ubK#j	  )��}�(h�K"j  ]�h�h�j  K#ubK$j	  )��}�(h�K"j  ]�h�h�j  K$ubK%j	  )��}�(h�K"j  ]�h�h�j  K%ubK&j	  )��}�(h�K"j  ]�h�h�j  K&ubK'j	  )��}�(h�K"j  ]�h�h�j  K'ubK(j	  )��}�(h�K"j  ]�h�h�j  K(ubK)j	  )��}�(h�K"j  ]�h�h�j  K)ubK*j	  )��}�(h�K"j  ]�h�h�j  K*ubK+j	  )��}�(h�K"j  ]�h�h�j  K+ubK,j	  )��}�(h�K"j  ]�h�h�j  K,ubK-j	  )��}�(h�K"j  ]�h�h�j  K-ubK.j	  )��}�(h�K"j  ]�h�h�j  K.ubK/j	  )��}�(h�K"j  ]�h�h�j  K/ubK0j	  )��}�(h�K"j  ]�h�h�j  K0ubK1j	  )��}�(h�K"j  ]�h�h�j  K1ubK2j	  )��}�(h�K"j  ]�h�h�j  K2ubK3j	  )��}�(h�K"j  ]�h�h�j  K3ubK4j	  )��}�(h�K"j  ]�h�h�j  K4ubK5j	  )��}�(h�K"j  ]�h�h�j  K5ubK6j	  )��}�(h�K"j  ]�h�h�j  K6ubK7j	  )��}�(h�K"j  ]�h�h�j  K7ubK8j	  )��}�(h�K"j  ]�h�h�j  K8ubK9j	  )��}�(h�K"j  ]�h�h�j  K9ubK:j	  )��}�(h�K"j  ]�h�h�j  K:ubK;j	  )��}�(h�K"j  ]�h�h�j  K;ubK<j	  )��}�(h�K"j  ]�h�h�j  K<ubK=j	  )��}�(h�K"j  ]�h�h�j  K=ubK>j	  )��}�(h�K"j  ]�h�h�j  K>ubK?j	  )��}�(h�K"j  ]�h�h�j  K?ubK@j	  )��}�(h�K"j  ]�h�h�j  K@ubKAj	  )��}�(h�K"j  ]�(KKeh�h�j  KAubKBj	  )��}�(h�K"j  ]�h�h�j  KBubKCj	  )��}�(h�K"j  ]�h�h�j  KCubuK#}�(K j	  )��}�(h�K#j  ]�h�h�j  K ubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubK	j	  )��}�(h�K#j  ]�h�h�j  K	ubK
j	  )��}�(h�K#j  ]�h�h�j  K
ubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubKj	  )��}�(h�K#j  ]�h�h�j  KubK j	  )��}�(h�K#j  ]�h�h�j  K ubK!j	  )��}�(h�K#j  ]�h�h�j  K!ubK"j	  )��}�(h�K#j  ]�h�h�j  K"ubK#j	  )��}�(h�K#j  ]�h�h�j  K#ubK$j	  )��}�(h�K#j  ]�h�h�j  K$ubK%j	  )��}�(h�K#j  ]�h�h�j  K%ubK&j	  )��}�(h�K#j  ]�h�h�j  K&ubK'j	  )��}�(h�K#j  ]�h�h�j  K'ubK(j	  )��}�(h�K#j  ]�h�h�j  K(ubK)j	  )��}�(h�K#j  ]�h�h�j  K)ubK*j	  )��}�(h�K#j  ]�h�h�j  K*ubK+j	  )��}�(h�K#j  ]�h�h�j  K+ubK,j	  )��}�(h�K#j  ]�h�h�j  K,ubK-j	  )��}�(h�K#j  ]�h�h�j  K-ubK.j	  )��}�(h�K#j  ]�h�h�j  K.ubK/j	  )��}�(h�K#j  ]�h�h�j  K/ubK0j	  )��}�(h�K#j  ]�h�h�j  K0ubK1j	  )��}�(h�K#j  ]�h�h�j  K1ubK2j	  )��}�(h�K#j  ]�h�h�j  K2ubK3j	  )��}�(h�K#j  ]�h�h�j  K3ubK4j	  )��}�(h�K#j  ]�h�h�j  K4ubK5j	  )��}�(h�K#j  ]�h�h�j  K5ubK6j	  )��}�(h�K#j  ]�h�h�j  K6ubK7j	  )��}�(h�K#j  ]�h�h�j  K7ubK8j	  )��}�(h�K#j  ]�h�h�j  K8ubK9j	  )��}�(h�K#j  ]�h�h�j  K9ubK:j	  )��}�(h�K#j  ]�h�h�j  K:ubK;j	  )��}�(h�K#j  ]�h�h�j  K;ubK<j	  )��}�(h�K#j  ]�h�h�j  K<ubK=j	  )��}�(h�K#j  ]�h�h�j  K=ubK>j	  )��}�(h�K#j  ]�h�h�j  K>ubK?j	  )��}�(h�K#j  ]�h�h�j  K?ubK@j	  )��}�(h�K#j  ]�h�h�j  K@ubKAj	  )��}�(h�K#j  ]�h�h�j  KAubKBj	  )��}�(h�K#j  ]�h�h�j  KBubKCj	  )��}�(h�K#j  ]�h�h�j  KCubuK$}�(K j	  )��}�(h�K$j  ]�h�h�j  K ubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubK	j	  )��}�(h�K$j  ]�h�h�j  K	ubK
j	  )��}�(h�K$j  ]�h�h�j  K
ubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubKj	  )��}�(h�K$j  ]�h�h�j  KubK j	  )��}�(h�K$j  ]�h�h�j  K ubK!j	  )��}�(h�K$j  ]�h�h�j  K!ubK"j	  )��}�(h�K$j  ]�h�h�j  K"ubK#j	  )��}�(h�K$j  ]�h�h�j  K#ubK$j	  )��}�(h�K$j  ]�h�h�j  K$ubK%j	  )��}�(h�K$j  ]�h�h�j  K%ubK&j	  )��}�(h�K$j  ]�h�h�j  K&ubK'j	  )��}�(h�K$j  ]�h�h�j  K'ubK(j	  )��}�(h�K$j  ]�h�h�j  K(ubK)j	  )��}�(h�K$j  ]�h�h�j  K)ubK*j	  )��}�(h�K$j  ]�h�h�j  K*ubK+j	  )��}�(h�K$j  ]�h�h�j  K+ubK,j	  )��}�(h�K$j  ]�h�h�j  K,ubK-j	  )��}�(h�K$j  ]�h�h�j  K-ubK.j	  )��}�(h�K$j  ]�h�h�j  K.ubK/j	  )��}�(h�K$j  ]�h�h�j  K/ubK0j	  )��}�(h�K$j  ]�h�h�j  K0ubK1j	  )��}�(h�K$j  ]�h�h�j  K1ubK2j	  )��}�(h�K$j  ]�h�h�j  K2ubK3j	  )��}�(h�K$j  ]�h�h�j  K3ubK4j	  )��}�(h�K$j  ]�h�h�j  K4ubK5j	  )��}�(h�K$j  ]�h�h�j  K5ubK6j	  )��}�(h�K$j  ]�h�h�j  K6ubK7j	  )��}�(h�K$j  ]�h�h�j  K7ubK8j	  )��}�(h�K$j  ]�h�h�j  K8ubK9j	  )��}�(h�K$j  ]�h�h�j  K9ubK:j	  )��}�(h�K$j  ]�h�h�j  K:ubK;j	  )��}�(h�K$j  ]�h�h�j  K;ubK<j	  )��}�(h�K$j  ]�h�h�j  K<ubK=j	  )��}�(h�K$j  ]�h�h�j  K=ubK>j	  )��}�(h�K$j  ]�h�h�j  K>ubK?j	  )��}�(h�K$j  ]�h�h�j  K?ubK@j	  )��}�(h�K$j  ]�h�h�j  K@ubKAj	  )��}�(h�K$j  ]�h�h�j  KAubKBj	  )��}�(h�K$j  ]�h�h�j  KBubKCj	  )��}�(h�K$j  ]�h�h�j  KCubuK%}�(K j	  )��}�(h�K%j  ]�h�h�j  K ubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubK	j	  )��}�(h�K%j  ]�h�h�j  K	ubK
j	  )��}�(h�K%j  ]�h�h�j  K
ubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubKj	  )��}�(h�K%j  ]�h�h�j  KubK j	  )��}�(h�K%j  ]�h�h�j  K ubK!j	  )��}�(h�K%j  ]�h�h�j  K!ubK"j	  )��}�(h�K%j  ]�h�h�j  K"ubK#j	  )��}�(h�K%j  ]�h�h�j  K#ubK$j	  )��}�(h�K%j  ]�h�h�j  K$ubK%j	  )��}�(h�K%j  ]�h�h�j  K%ubK&j	  )��}�(h�K%j  ]�h�h�j  K&ubK'j	  )��}�(h�K%j  ]�h�h�j  K'ubK(j	  )��}�(h�K%j  ]�h�h�j  K(ubK)j	  )��}�(h�K%j  ]�h�h�j  K)ubK*j	  )��}�(h�K%j  ]�h�h�j  K*ubK+j	  )��}�(h�K%j  ]�h�h�j  K+ubK,j	  )��}�(h�K%j  ]�h�h�j  K,ubK-j	  )��}�(h�K%j  ]�h�h�j  K-ubK.j	  )��}�(h�K%j  ]�h�h�j  K.ubK/j	  )��}�(h�K%j  ]�h�h�j  K/ubK0j	  )��}�(h�K%j  ]�h�h�j  K0ubK1j	  )��}�(h�K%j  ]�h�h�j  K1ubK2j	  )��}�(h�K%j  ]�h�h�j  K2ubK3j	  )��}�(h�K%j  ]�h�h�j  K3ubK4j	  )��}�(h�K%j  ]�h�h�j  K4ubK5j	  )��}�(h�K%j  ]�h�h�j  K5ubK6j	  )��}�(h�K%j  ]�h�h�j  K6ubK7j	  )��}�(h�K%j  ]�h�h�j  K7ubK8j	  )��}�(h�K%j  ]�h�h�j  K8ubK9j	  )��}�(h�K%j  ]�h�h�j  K9ubK:j	  )��}�(h�K%j  ]�h�h�j  K:ubK;j	  )��}�(h�K%j  ]�h�h�j  K;ubK<j	  )��}�(h�K%j  ]�h�h�j  K<ubK=j	  )��}�(h�K%j  ]�h�h�j  K=ubK>j	  )��}�(h�K%j  ]�h�h�j  K>ubK?j	  )��}�(h�K%j  ]�h�h�j  K?ubK@j	  )��}�(h�K%j  ]�h�h�j  K@ubKAj	  )��}�(h�K%j  ]�h�h�j  KAubKBj	  )��}�(h�K%j  ]�h�h�j  KBubKCj	  )��}�(h�K%j  ]�h�h�j  KCubuK&}�(K j	  )��}�(h�K&j  ]�h�h�j  K ubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubK	j	  )��}�(h�K&j  ]�h�h�j  K	ubK
j	  )��}�(h�K&j  ]�h�h�j  K
ubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubKj	  )��}�(h�K&j  ]�h�h�j  KubK j	  )��}�(h�K&j  ]�h�h�j  K ubK!j	  )��}�(h�K&j  ]�h�h�j  K!ubK"j	  )��}�(h�K&j  ]�h�h�j  K"ubK#j	  )��}�(h�K&j  ]�h�h�j  K#ubK$j	  )��}�(h�K&j  ]�h�h�j  K$ubK%j	  )��}�(h�K&j  ]�h�h�j  K%ubK&j	  )��}�(h�K&j  ]�h�h�j  K&ubK'j	  )��}�(h�K&j  ]�h�h�j  K'ubK(j	  )��}�(h�K&j  ]�h�h�j  K(ubK)j	  )��}�(h�K&j  ]�h�h�j  K)ubK*j	  )��}�(h�K&j  ]�h�h�j  K*ubK+j	  )��}�(h�K&j  ]�h�h�j  K+ubK,j	  )��}�(h�K&j  ]�h�h�j  K,ubK-j	  )��}�(h�K&j  ]�h�h�j  K-ubK.j	  )��}�(h�K&j  ]�h�h�j  K.ubK/j	  )��}�(h�K&j  ]�h�h�j  K/ubK0j	  )��}�(h�K&j  ]�h�h�j  K0ubK1j	  )��}�(h�K&j  ]�h�h�j  K1ubK2j	  )��}�(h�K&j  ]�h�h�j  K2ubK3j	  )��}�(h�K&j  ]�h�h�j  K3ubK4j	  )��}�(h�K&j  ]�h�h�j  K4ubK5j	  )��}�(h�K&j  ]�h�h�j  K5ubK6j	  )��}�(h�K&j  ]�h�h�j  K6ubK7j	  )��}�(h�K&j  ]�h�h�j  K7ubK8j	  )��}�(h�K&j  ]�h�h�j  K8ubK9j	  )��}�(h�K&j  ]�h�h�j  K9ubK:j	  )��}�(h�K&j  ]�h�h�j  K:ubK;j	  )��}�(h�K&j  ]�h�h�j  K;ubK<j	  )��}�(h�K&j  ]�h�h�j  K<ubK=j	  )��}�(h�K&j  ]�h�h�j  K=ubK>j	  )��}�(h�K&j  ]�h�h�j  K>ubK?j	  )��}�(h�K&j  ]�h�h�j  K?ubK@j	  )��}�(h�K&j  ]�h�h�j  K@ubKAj	  )��}�(h�K&j  ]�h�h�j  KAubKBj	  )��}�(h�K&j  ]�h�h�j  KBubKCj	  )��}�(h�K&j  ]�h�h�j  KCubuK'}�(K j	  )��}�(h�K'j  ]�h�h�j  K ubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubK	j	  )��}�(h�K'j  ]�h�h�j  K	ubK
j	  )��}�(h�K'j  ]�h�h�j  K
ubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubKj	  )��}�(h�K'j  ]�h�h�j  KubK j	  )��}�(h�K'j  ]�h�h�j  K ubK!j	  )��}�(h�K'j  ]�h�h�j  K!ubK"j	  )��}�(h�K'j  ]�h�h�j  K"ubK#j	  )��}�(h�K'j  ]�h�h�j  K#ubK$j	  )��}�(h�K'j  ]�h�h�j  K$ubK%j	  )��}�(h�K'j  ]�h�h�j  K%ubK&j	  )��}�(h�K'j  ]�h�h�j  K&ubK'j	  )��}�(h�K'j  ]�h�h�j  K'ubK(j	  )��}�(h�K'j  ]�h�h�j  K(ubK)j	  )��}�(h�K'j  ]�h�h�j  K)ubK*j	  )��}�(h�K'j  ]�h�h�j  K*ubK+j	  )��}�(h�K'j  ]�h�h�j  K+ubK,j	  )��}�(h�K'j  ]�h�h�j  K,ubK-j	  )��}�(h�K'j  ]�h�h�j  K-ubK.j	  )��}�(h�K'j  ]�h�h�j  K.ubK/j	  )��}�(h�K'j  ]�h�h�j  K/ubK0j	  )��}�(h�K'j  ]�h�h�j  K0ubK1j	  )��}�(h�K'j  ]�h�h�j  K1ubK2j	  )��}�(h�K'j  ]�h�h�j  K2ubK3j	  )��}�(h�K'j  ]�h�h�j  K3ubK4j	  )��}�(h�K'j  ]�h�h�j  K4ubK5j	  )��}�(h�K'j  ]�h�h�j  K5ubK6j	  )��}�(h�K'j  ]�h�h�j  K6ubK7j	  )��}�(h�K'j  ]�h�h�j  K7ubK8j	  )��}�(h�K'j  ]�h�h�j  K8ubK9j	  )��}�(h�K'j  ]�h�h�j  K9ubK:j	  )��}�(h�K'j  ]�h�h�j  K:ubK;j	  )��}�(h�K'j  ]�h�h�j  K;ubK<j	  )��}�(h�K'j  ]�h�h�j  K<ubK=j	  )��}�(h�K'j  ]�h�h�j  K=ubK>j	  )��}�(h�K'j  ]�h�h�j  K>ubK?j	  )��}�(h�K'j  ]�h�h�j  K?ubK@j	  )��}�(h�K'j  ]�h�h�j  K@ubKAj	  )��}�(h�K'j  ]�h�h�j  KAubKBj	  )��}�(h�K'j  ]�h�h�j  KBubKCj	  )��}�(h�K'j  ]�h�h�j  KCubuK(}�(K j	  )��}�(h�K(j  ]�h�h�j  K ubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubK	j	  )��}�(h�K(j  ]�h�h�j  K	ubK
j	  )��}�(h�K(j  ]�h�h�j  K
ubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubKj	  )��}�(h�K(j  ]�h�h�j  KubK j	  )��}�(h�K(j  ]�h�h�j  K ubK!j	  )��}�(h�K(j  ]�h�h�j  K!ubK"j	  )��}�(h�K(j  ]�h�h�j  K"ubK#j	  )��}�(h�K(j  ]�h�h�j  K#ubK$j	  )��}�(h�K(j  ]�h�h�j  K$ubK%j	  )��}�(h�K(j  ]�h�h�j  K%ubK&j	  )��}�(h�K(j  ]�h�h�j  K&ubK'j	  )��}�(h�K(j  ]�h�h�j  K'ubK(j	  )��}�(h�K(j  ]�h�h�j  K(ubK)j	  )��}�(h�K(j  ]�h�h�j  K)ubK*j	  )��}�(h�K(j  ]�h�h�j  K*ubK+j	  )��}�(h�K(j  ]�h�h�j  K+ubK,j	  )��}�(h�K(j  ]�h�h�j  K,ubK-j	  )��}�(h�K(j  ]�h�h�j  K-ubK.j	  )��}�(h�K(j  ]�h�h�j  K.ubK/j	  )��}�(h�K(j  ]�h�h�j  K/ubK0j	  )��}�(h�K(j  ]�h�h�j  K0ubK1j	  )��}�(h�K(j  ]�h�h�j  K1ubK2j	  )��}�(h�K(j  ]�h�h�j  K2ubK3j	  )��}�(h�K(j  ]�h�h�j  K3ubK4j	  )��}�(h�K(j  ]�h�h�j  K4ubK5j	  )��}�(h�K(j  ]�h�h�j  K5ubK6j	  )��}�(h�K(j  ]�h�h�j  K6ubK7j	  )��}�(h�K(j  ]�h�h�j  K7ubK8j	  )��}�(h�K(j  ]�h�h�j  K8ubK9j	  )��}�(h�K(j  ]�h�h�j  K9ubK:j	  )��}�(h�K(j  ]�h�h�j  K:ubK;j	  )��}�(h�K(j  ]�h�h�j  K;ubK<j	  )��}�(h�K(j  ]�h�h�j  K<ubK=j	  )��}�(h�K(j  ]�h�h�j  K=ubK>j	  )��}�(h�K(j  ]�h�h�j  K>ubK?j	  )��}�(h�K(j  ]�h�h�j  K?ubK@j	  )��}�(h�K(j  ]�h�h�j  K@ubKAj	  )��}�(h�K(j  ]�h�h�j  KAubKBj	  )��}�(h�K(j  ]�h�h�j  KBubKCj	  )��}�(h�K(j  ]�h�h�j  KCubuK)}�(K j	  )��}�(h�K)j  ]�h�h�j  K ubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubK	j	  )��}�(h�K)j  ]�h�h�j  K	ubK
j	  )��}�(h�K)j  ]�h�h�j  K
ubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubKj	  )��}�(h�K)j  ]�h�h�j  KubK j	  )��}�(h�K)j  ]�h�h�j  K ubK!j	  )��}�(h�K)j  ]�h�h�j  K!ubK"j	  )��}�(h�K)j  ]�h�h�j  K"ubK#j	  )��}�(h�K)j  ]�h�h�j  K#ubK$j	  )��}�(h�K)j  ]�h�h�j  K$ubK%j	  )��}�(h�K)j  ]�h�h�j  K%ubK&j	  )��}�(h�K)j  ]�h�h�j  K&ubK'j	  )��}�(h�K)j  ]�h�h�j  K'ubK(j	  )��}�(h�K)j  ]�h�h�j  K(ubK)j	  )��}�(h�K)j  ]�h�h�j  K)ubK*j	  )��}�(h�K)j  ]�h�h�j  K*ubK+j	  )��}�(h�K)j  ]�h�h�j  K+ubK,j	  )��}�(h�K)j  ]�h�h�j  K,ubK-j	  )��}�(h�K)j  ]�h�h�j  K-ubK.j	  )��}�(h�K)j  ]�h�h�j  K.ubK/j	  )��}�(h�K)j  ]�h�h�j  K/ubK0j	  )��}�(h�K)j  ]�h�h�j  K0ubK1j	  )��}�(h�K)j  ]�h�h�j  K1ubK2j	  )��}�(h�K)j  ]�h�h�j  K2ubK3j	  )��}�(h�K)j  ]�h�h�j  K3ubK4j	  )��}�(h�K)j  ]�h�h�j  K4ubK5j	  )��}�(h�K)j  ]�h�h�j  K5ubK6j	  )��}�(h�K)j  ]�h�h�j  K6ubK7j	  )��}�(h�K)j  ]�h�h�j  K7ubK8j	  )��}�(h�K)j  ]�h�h�j  K8ubK9j	  )��}�(h�K)j  ]�h�h�j  K9ubK:j	  )��}�(h�K)j  ]�h�h�j  K:ubK;j	  )��}�(h�K)j  ]�h�h�j  K;ubK<j	  )��}�(h�K)j  ]�h�h�j  K<ubK=j	  )��}�(h�K)j  ]�h�h�j  K=ubK>j	  )��}�(h�K)j  ]�h�h�j  K>ubK?j	  )��}�(h�K)j  ]�h�h�j  K?ubK@j	  )��}�(h�K)j  ]�h�h�j  K@ubKAj	  )��}�(h�K)j  ]�h�h�j  KAubKBj	  )��}�(h�K)j  ]�h�h�j  KBubKCj	  )��}�(h�K)j  ]�h�h�j  KCubuK*}�(K j	  )��}�(h�K*j  ]�h�h�j  K ubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubK	j	  )��}�(h�K*j  ]�h�h�j  K	ubK
j	  )��}�(h�K*j  ]�h�h�j  K
ubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubKj	  )��}�(h�K*j  ]�h�h�j  KubK j	  )��}�(h�K*j  ]�h�h�j  K ubK!j	  )��}�(h�K*j  ]�h�h�j  K!ubK"j	  )��}�(h�K*j  ]�h�h�j  K"ubK#j	  )��}�(h�K*j  ]�h�h�j  K#ubK$j	  )��}�(h�K*j  ]�h�h�j  K$ubK%j	  )��}�(h�K*j  ]�h�h�j  K%ubK&j	  )��}�(h�K*j  ]�h�h�j  K&ubK'j	  )��}�(h�K*j  ]�h�h�j  K'ubK(j	  )��}�(h�K*j  ]�h�h�j  K(ubK)j	  )��}�(h�K*j  ]�h�h�j  K)ubK*j	  )��}�(h�K*j  ]�h�h�j  K*ubK+j	  )��}�(h�K*j  ]�h�h�j  K+ubK,j	  )��}�(h�K*j  ]�h�h�j  K,ubK-j	  )��}�(h�K*j  ]�h�h�j  K-ubK.j	  )��}�(h�K*j  ]�h�h�j  K.ubK/j	  )��}�(h�K*j  ]�h�h�j  K/ubK0j	  )��}�(h�K*j  ]�h�h�j  K0ubK1j	  )��}�(h�K*j  ]�h�h�j  K1ubK2j	  )��}�(h�K*j  ]�h�h�j  K2ubK3j	  )��}�(h�K*j  ]�h�h�j  K3ubK4j	  )��}�(h�K*j  ]�h�h�j  K4ubK5j	  )��}�(h�K*j  ]�h�h�j  K5ubK6j	  )��}�(h�K*j  ]�h�h�j  K6ubK7j	  )��}�(h�K*j  ]�h�h�j  K7ubK8j	  )��}�(h�K*j  ]�h�h�j  K8ubK9j	  )��}�(h�K*j  ]�h�h�j  K9ubK:j	  )��}�(h�K*j  ]�h�h�j  K:ubK;j	  )��}�(h�K*j  ]�h�h�j  K;ubK<j	  )��}�(h�K*j  ]�h�h�j  K<ubK=j	  )��}�(h�K*j  ]�h�h�j  K=ubK>j	  )��}�(h�K*j  ]�h�h�j  K>ubK?j	  )��}�(h�K*j  ]�h�h�j  K?ubK@j	  )��}�(h�K*j  ]�h�h�j  K@ubKAj	  )��}�(h�K*j  ]�h�h�j  KAubKBj	  )��}�(h�K*j  ]�h�h�j  KBubKCj	  )��}�(h�K*j  ]�h�h�j  KCubuK+}�(K j	  )��}�(h�K+j  ]�h�h�j  K ubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubK	j	  )��}�(h�K+j  ]�h�h�j  K	ubK
j	  )��}�(h�K+j  ]�h�h�j  K
ubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubKj	  )��}�(h�K+j  ]�h�h�j  KubK j	  )��}�(h�K+j  ]�h�h�j  K ubK!j	  )��}�(h�K+j  ]�h�h�j  K!ubK"j	  )��}�(h�K+j  ]�h�h�j  K"ubK#j	  )��}�(h�K+j  ]�h�h�j  K#ubK$j	  )��}�(h�K+j  ]�h�h�j  K$ubK%j	  )��}�(h�K+j  ]�h�h�j  K%ubK&j	  )��}�(h�K+j  ]�h�h�j  K&ubK'j	  )��}�(h�K+j  ]�h�h�j  K'ubK(j	  )��}�(h�K+j  ]�h�h�j  K(ubK)j	  )��}�(h�K+j  ]�h�h�j  K)ubK*j	  )��}�(h�K+j  ]�h�h�j  K*ubK+j	  )��}�(h�K+j  ]�h�h�j  K+ubK,j	  )��}�(h�K+j  ]�h�h�j  K,ubK-j	  )��}�(h�K+j  ]�h�h�j  K-ubK.j	  )��}�(h�K+j  ]�h�h�j  K.ubK/j	  )��}�(h�K+j  ]�h�h�j  K/ubK0j	  )��}�(h�K+j  ]�h�h�j  K0ubK1j	  )��}�(h�K+j  ]�h�h�j  K1ubK2j	  )��}�(h�K+j  ]�h�h�j  K2ubK3j	  )��}�(h�K+j  ]�h�h�j  K3ubK4j	  )��}�(h�K+j  ]�h�h�j  K4ubK5j	  )��}�(h�K+j  ]�h�h�j  K5ubK6j	  )��}�(h�K+j  ]�h�h�j  K6ubK7j	  )��}�(h�K+j  ]�h�h�j  K7ubK8j	  )��}�(h�K+j  ]�h�h�j  K8ubK9j	  )��}�(h�K+j  ]�h�h�j  K9ubK:j	  )��}�(h�K+j  ]�h�h�j  K:ubK;j	  )��}�(h�K+j  ]�h�h�j  K;ubK<j	  )��}�(h�K+j  ]�h�h�j  K<ubK=j	  )��}�(h�K+j  ]�h�h�j  K=ubK>j	  )��}�(h�K+j  ]�h�h�j  K>ubK?j	  )��}�(h�K+j  ]�h�h�j  K?ubK@j	  )��}�(h�K+j  ]�h�h�j  K@ubKAj	  )��}�(h�K+j  ]�h�h�j  KAubKBj	  )��}�(h�K+j  ]�h�h�j  KBubKCj	  )��}�(h�K+j  ]�h�h�j  KCubuK,}�(K j	  )��}�(h�K,j  ]�h�h�j  K ubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubK	j	  )��}�(h�K,j  ]�h�h�j  K	ubK
j	  )��}�(h�K,j  ]�h�h�j  K
ubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubKj	  )��}�(h�K,j  ]�h�h�j  KubK j	  )��}�(h�K,j  ]�h�h�j  K ubK!j	  )��}�(h�K,j  ]�h�h�j  K!ubK"j	  )��}�(h�K,j  ]�h�h�j  K"ubK#j	  )��}�(h�K,j  ]�h�h�j  K#ubK$j	  )��}�(h�K,j  ]�h�h�j  K$ubK%j	  )��}�(h�K,j  ]�h�h�j  K%ubK&j	  )��}�(h�K,j  ]�h�h�j  K&ubK'j	  )��}�(h�K,j  ]�h�h�j  K'ubK(j	  )��}�(h�K,j  ]�h�h�j  K(ubK)j	  )��}�(h�K,j  ]�h�h�j  K)ubK*j	  )��}�(h�K,j  ]�h�h�j  K*ubK+j	  )��}�(h�K,j  ]�h�h�j  K+ubK,j	  )��}�(h�K,j  ]�h�h�j  K,ubK-j	  )��}�(h�K,j  ]�h�h�j  K-ubK.j	  )��}�(h�K,j  ]�h�h�j  K.ubK/j	  )��}�(h�K,j  ]�h�h�j  K/ubK0j	  )��}�(h�K,j  ]�h�h�j  K0ubK1j	  )��}�(h�K,j  ]�h�h�j  K1ubK2j	  )��}�(h�K,j  ]�h�h�j  K2ubK3j	  )��}�(h�K,j  ]�h�h�j  K3ubK4j	  )��}�(h�K,j  ]�h�h�j  K4ubK5j	  )��}�(h�K,j  ]�h�h�j  K5ubK6j	  )��}�(h�K,j  ]�h�h�j  K6ubK7j	  )��}�(h�K,j  ]�h�h�j  K7ubK8j	  )��}�(h�K,j  ]�h�h�j  K8ubK9j	  )��}�(h�K,j  ]�h�h�j  K9ubK:j	  )��}�(h�K,j  ]�h�h�j  K:ubK;j	  )��}�(h�K,j  ]�h�h�j  K;ubK<j	  )��}�(h�K,j  ]�h�h�j  K<ubK=j	  )��}�(h�K,j  ]�h�h�j  K=ubK>j	  )��}�(h�K,j  ]�h�h�j  K>ubK?j	  )��}�(h�K,j  ]�h�h�j  K?ubK@j	  )��}�(h�K,j  ]�h�h�j  K@ubKAj	  )��}�(h�K,j  ]�h�h�j  KAubKBj	  )��}�(h�K,j  ]�h�h�j  KBubKCj	  )��}�(h�K,j  ]�h�h�j  KCubuK-}�(K j	  )��}�(h�K-j  ]�h�h�j  K ubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubK	j	  )��}�(h�K-j  ]�h�h�j  K	ubK
j	  )��}�(h�K-j  ]�h�h�j  K
ubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubKj	  )��}�(h�K-j  ]�h�h�j  KubK j	  )��}�(h�K-j  ]�h�h�j  K ubK!j	  )��}�(h�K-j  ]�h�h�j  K!ubK"j	  )��}�(h�K-j  ]�h�h�j  K"ubK#j	  )��}�(h�K-j  ]�h�h�j  K#ubK$j	  )��}�(h�K-j  ]�h�h�j  K$ubK%j	  )��}�(h�K-j  ]�h�h�j  K%ubK&j	  )��}�(h�K-j  ]�h�h�j  K&ubK'j	  )��}�(h�K-j  ]�h�h�j  K'ubK(j	  )��}�(h�K-j  ]�h�h�j  K(ubK)j	  )��}�(h�K-j  ]�h�h�j  K)ubK*j	  )��}�(h�K-j  ]�h�h�j  K*ubK+j	  )��}�(h�K-j  ]�h�h�j  K+ubK,j	  )��}�(h�K-j  ]�h�h�j  K,ubK-j	  )��}�(h�K-j  ]�h�h�j  K-ubK.j	  )��}�(h�K-j  ]�h�h�j  K.ubK/j	  )��}�(h�K-j  ]�h�h�j  K/ubK0j	  )��}�(h�K-j  ]�h�h�j  K0ubK1j	  )��}�(h�K-j  ]�h�h�j  K1ubK2j	  )��}�(h�K-j  ]�h�h�j  K2ubK3j	  )��}�(h�K-j  ]�h�h�j  K3ubK4j	  )��}�(h�K-j  ]�h�h�j  K4ubK5j	  )��}�(h�K-j  ]�h�h�j  K5ubK6j	  )��}�(h�K-j  ]�h�h�j  K6ubK7j	  )��}�(h�K-j  ]�h�h�j  K7ubK8j	  )��}�(h�K-j  ]�h�h�j  K8ubK9j	  )��}�(h�K-j  ]�h�h�j  K9ubK:j	  )��}�(h�K-j  ]�h�h�j  K:ubK;j	  )��}�(h�K-j  ]�h�h�j  K;ubK<j	  )��}�(h�K-j  ]�h�h�j  K<ubK=j	  )��}�(h�K-j  ]�h�h�j  K=ubK>j	  )��}�(h�K-j  ]�h�h�j  K>ubK?j	  )��}�(h�K-j  ]�h�h�j  K?ubK@j	  )��}�(h�K-j  ]�h�h�j  K@ubKAj	  )��}�(h�K-j  ]�h�h�j  KAubKBj	  )��}�(h�K-j  ]�h�h�j  KBubKCj	  )��}�(h�K-j  ]�h�h�j  KCubuK.}�(K j	  )��}�(h�K.j  ]�h�h�j  K ubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubK	j	  )��}�(h�K.j  ]�h�h�j  K	ubK
j	  )��}�(h�K.j  ]�h�h�j  K
ubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubKj	  )��}�(h�K.j  ]�h�h�j  KubK j	  )��}�(h�K.j  ]�h�h�j  K ubK!j	  )��}�(h�K.j  ]�h�h�j  K!ubK"j	  )��}�(h�K.j  ]�h�h�j  K"ubK#j	  )��}�(h�K.j  ]�h�h�j  K#ubK$j	  )��}�(h�K.j  ]�h�h�j  K$ubK%j	  )��}�(h�K.j  ]�h�h�j  K%ubK&j	  )��}�(h�K.j  ]�h�h�j  K&ubK'j	  )��}�(h�K.j  ]�h�h�j  K'ubK(j	  )��}�(h�K.j  ]�h�h�j  K(ubK)j	  )��}�(h�K.j  ]�h�h�j  K)ubK*j	  )��}�(h�K.j  ]�h�h�j  K*ubK+j	  )��}�(h�K.j  ]�h�h�j  K+ubK,j	  )��}�(h�K.j  ]�h�h�j  K,ubK-j	  )��}�(h�K.j  ]�h�h�j  K-ubK.j	  )��}�(h�K.j  ]�h�h�j  K.ubK/j	  )��}�(h�K.j  ]�h�h�j  K/ubK0j	  )��}�(h�K.j  ]�h�h�j  K0ubK1j	  )��}�(h�K.j  ]�h�h�j  K1ubK2j	  )��}�(h�K.j  ]�h�h�j  K2ubK3j	  )��}�(h�K.j  ]�h�h�j  K3ubK4j	  )��}�(h�K.j  ]�h�h�j  K4ubK5j	  )��}�(h�K.j  ]�h�h�j  K5ubK6j	  )��}�(h�K.j  ]�h�h�j  K6ubK7j	  )��}�(h�K.j  ]�h�h�j  K7ubK8j	  )��}�(h�K.j  ]�h�h�j  K8ubK9j	  )��}�(h�K.j  ]�h�h�j  K9ubK:j	  )��}�(h�K.j  ]�h�h�j  K:ubK;j	  )��}�(h�K.j  ]�h�h�j  K;ubK<j	  )��}�(h�K.j  ]�h�h�j  K<ubK=j	  )��}�(h�K.j  ]�h�h�j  K=ubK>j	  )��}�(h�K.j  ]�h�h�j  K>ubK?j	  )��}�(h�K.j  ]�h�h�j  K?ubK@j	  )��}�(h�K.j  ]�h�h�j  K@ubKAj	  )��}�(h�K.j  ]�h�h�j  KAubKBj	  )��}�(h�K.j  ]�h�h�j  KBubKCj	  )��}�(h�K.j  ]�h�h�j  KCubuK/}�(K j	  )��}�(h�K/j  ]�h�h�j  K ubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubK	j	  )��}�(h�K/j  ]�h�h�j  K	ubK
j	  )��}�(h�K/j  ]�h�h�j  K
ubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubKj	  )��}�(h�K/j  ]�h�h�j  KubK j	  )��}�(h�K/j  ]�h�h�j  K ubK!j	  )��}�(h�K/j  ]�h�h�j  K!ubK"j	  )��}�(h�K/j  ]�h�h�j  K"ubK#j	  )��}�(h�K/j  ]�h�h�j  K#ubK$j	  )��}�(h�K/j  ]�h�h�j  K$ubK%j	  )��}�(h�K/j  ]�h�h�j  K%ubK&j	  )��}�(h�K/j  ]�h�h�j  K&ubK'j	  )��}�(h�K/j  ]�h�h�j  K'ubK(j	  )��}�(h�K/j  ]�h�h�j  K(ubK)j	  )��}�(h�K/j  ]�h�h�j  K)ubK*j	  )��}�(h�K/j  ]�h�h�j  K*ubK+j	  )��}�(h�K/j  ]�h�h�j  K+ubK,j	  )��}�(h�K/j  ]�h�h�j  K,ubK-j	  )��}�(h�K/j  ]�h�h�j  K-ubK.j	  )��}�(h�K/j  ]�h�h�j  K.ubK/j	  )��}�(h�K/j  ]�h�h�j  K/ubK0j	  )��}�(h�K/j  ]�h�h�j  K0ubK1j	  )��}�(h�K/j  ]�h�h�j  K1ubK2j	  )��}�(h�K/j  ]�h�h�j  K2ubK3j	  )��}�(h�K/j  ]�h�h�j  K3ubK4j	  )��}�(h�K/j  ]�h�h�j  K4ubK5j	  )��}�(h�K/j  ]�h�h�j  K5ubK6j	  )��}�(h�K/j  ]�h�h�j  K6ubK7j	  )��}�(h�K/j  ]�h�h�j  K7ubK8j	  )��}�(h�K/j  ]�h�h�j  K8ubK9j	  )��}�(h�K/j  ]�h�h�j  K9ubK:j	  )��}�(h�K/j  ]�h�h�j  K:ubK;j	  )��}�(h�K/j  ]�h�h�j  K;ubK<j	  )��}�(h�K/j  ]�h�h�j  K<ubK=j	  )��}�(h�K/j  ]�h�h�j  K=ubK>j	  )��}�(h�K/j  ]�h�h�j  K>ubK?j	  )��}�(h�K/j  ]�h�h�j  K?ubK@j	  )��}�(h�K/j  ]�h�h�j  K@ubKAj	  )��}�(h�K/j  ]�h�h�j  KAubKBj	  )��}�(h�K/j  ]�h�h�j  KBubKCj	  )��}�(h�K/j  ]�h�h�j  KCubuK0}�(K j	  )��}�(h�K0j  ]�h�h�j  K ubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubK	j	  )��}�(h�K0j  ]�h�h�j  K	ubK
j	  )��}�(h�K0j  ]�h�h�j  K
ubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubKj	  )��}�(h�K0j  ]�h�h�j  KubK j	  )��}�(h�K0j  ]�h�h�j  K ubK!j	  )��}�(h�K0j  ]�h�h�j  K!ubK"j	  )��}�(h�K0j  ]�h�h�j  K"ubK#j	  )��}�(h�K0j  ]�h�h�j  K#ubK$j	  )��}�(h�K0j  ]�h�h�j  K$ubK%j	  )��}�(h�K0j  ]�h�h�j  K%ubK&j	  )��}�(h�K0j  ]�h�h�j  K&ubK'j	  )��}�(h�K0j  ]�h�h�j  K'ubK(j	  )��}�(h�K0j  ]�h�h�j  K(ubK)j	  )��}�(h�K0j  ]�h�h�j  K)ubK*j	  )��}�(h�K0j  ]�h�h�j  K*ubK+j	  )��}�(h�K0j  ]�h�h�j  K+ubK,j	  )��}�(h�K0j  ]�h�h�j  K,ubK-j	  )��}�(h�K0j  ]�h�h�j  K-ubK.j	  )��}�(h�K0j  ]�h�h�j  K.ubK/j	  )��}�(h�K0j  ]�h�h�j  K/ubK0j	  )��}�(h�K0j  ]�h�h�j  K0ubK1j	  )��}�(h�K0j  ]�h�h�j  K1ubK2j	  )��}�(h�K0j  ]�h�h�j  K2ubK3j	  )��}�(h�K0j  ]�h�h�j  K3ubK4j	  )��}�(h�K0j  ]�h�h�j  K4ubK5j	  )��}�(h�K0j  ]�h�h�j  K5ubK6j	  )��}�(h�K0j  ]�h�h�j  K6ubK7j	  )��}�(h�K0j  ]�h�h�j  K7ubK8j	  )��}�(h�K0j  ]�h�h�j  K8ubK9j	  )��}�(h�K0j  ]�h�h�j  K9ubK:j	  )��}�(h�K0j  ]�h�h�j  K:ubK;j	  )��}�(h�K0j  ]�h�h�j  K;ubK<j	  )��}�(h�K0j  ]�h�h�j  K<ubK=j	  )��}�(h�K0j  ]�h�h�j  K=ubK>j	  )��}�(h�K0j  ]�h�h�j  K>ubK?j	  )��}�(h�K0j  ]�h�h�j  K?ubK@j	  )��}�(h�K0j  ]�h�h�j  K@ubKAj	  )��}�(h�K0j  ]�h�h�j  KAubKBj	  )��}�(h�K0j  ]�h�h�j  KBubKCj	  )��}�(h�K0j  ]�h�h�j  KCubuK1}�(K j	  )��}�(h�K1j  ]�h�h�j  K ubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubK	j	  )��}�(h�K1j  ]�h�h�j  K	ubK
j	  )��}�(h�K1j  ]�h�h�j  K
ubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubKj	  )��}�(h�K1j  ]�h�h�j  KubK j	  )��}�(h�K1j  ]�h�h�j  K ubK!j	  )��}�(h�K1j  ]�h�h�j  K!ubK"j	  )��}�(h�K1j  ]�h�h�j  K"ubK#j	  )��}�(h�K1j  ]�h�h�j  K#ubK$j	  )��}�(h�K1j  ]�h�h�j  K$ubK%j	  )��}�(h�K1j  ]�h�h�j  K%ubK&j	  )��}�(h�K1j  ]�h�h�j  K&ubK'j	  )��}�(h�K1j  ]�h�h�j  K'ubK(j	  )��}�(h�K1j  ]�h�h�j  K(ubK)j	  )��}�(h�K1j  ]�h�h�j  K)ubK*j	  )��}�(h�K1j  ]�h�h�j  K*ubK+j	  )��}�(h�K1j  ]�h�h�j  K+ubK,j	  )��}�(h�K1j  ]�h�h�j  K,ubK-j	  )��}�(h�K1j  ]�h�h�j  K-ubK.j	  )��}�(h�K1j  ]�h�h�j  K.ubK/j	  )��}�(h�K1j  ]�h�h�j  K/ubK0j	  )��}�(h�K1j  ]�h�h�j  K0ubK1j	  )��}�(h�K1j  ]�h�h�j  K1ubK2j	  )��}�(h�K1j  ]�h�h�j  K2ubK3j	  )��}�(h�K1j  ]�h�h�j  K3ubK4j	  )��}�(h�K1j  ]�h�h�j  K4ubK5j	  )��}�(h�K1j  ]�h�h�j  K5ubK6j	  )��}�(h�K1j  ]�h�h�j  K6ubK7j	  )��}�(h�K1j  ]�h�h�j  K7ubK8j	  )��}�(h�K1j  ]�h�h�j  K8ubK9j	  )��}�(h�K1j  ]�h�h�j  K9ubK:j	  )��}�(h�K1j  ]�h�h�j  K:ubK;j	  )��}�(h�K1j  ]�h�h�j  K;ubK<j	  )��}�(h�K1j  ]�h�h�j  K<ubK=j	  )��}�(h�K1j  ]�h�h�j  K=ubK>j	  )��}�(h�K1j  ]�h�h�j  K>ubK?j	  )��}�(h�K1j  ]�h�h�j  K?ubK@j	  )��}�(h�K1j  ]�h�h�j  K@ubKAj	  )��}�(h�K1j  ]�h�h�j  KAubKBj	  )��}�(h�K1j  ]�h�h�j  KBubKCj	  )��}�(h�K1j  ]�h�h�j  KCubuK2}�(K j	  )��}�(h�K2j  ]�h�h�j  K ubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubK	j	  )��}�(h�K2j  ]�h�h�j  K	ubK
j	  )��}�(h�K2j  ]�h�h�j  K
ubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )���       }�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubKj	  )��}�(h�K2j  ]�h�h�j  KubK j	  )��}�(h�K2j  ]�h�h�j  K ubK!j	  )��}�(h�K2j  ]�h�h�j  K!ubK"j	  )��}�(h�K2j  ]�h�h�j  K"ubK#j	  )��}�(h�K2j  ]�h�h�j  K#ubK$j	  )��}�(h�K2j  ]�h�h�j  K$ubK%j	  )��}�(h�K2j  ]�h�h�j  K%ubK&j	  )��}�(h�K2j  ]�h�h�j  K&ubK'j	  )��}�(h�K2j  ]�h�h�j  K'ubK(j	  )��}�(h�K2j  ]�h�h�j  K(ubK)j	  )��}�(h�K2j  ]�h�h�j  K)ubK*j	  )��}�(h�K2j  ]�h�h�j  K*ubK+j	  )��}�(h�K2j  ]�h�h�j  K+ubK,j	  )��}�(h�K2j  ]�h�h�j  K,ubK-j	  )��}�(h�K2j  ]�h�h�j  K-ubK.j	  )��}�(h�K2j  ]�h�h�j  K.ubK/j	  )��}�(h�K2j  ]�h�h�j  K/ubK0j	  )��}�(h�K2j  ]�h�h�j  K0ubK1j	  )��}�(h�K2j  ]�h�h�j  K1ubK2j	  )��}�(h�K2j  ]�h�h�j  K2ubK3j	  )��}�(h�K2j  ]�h�h�j  K3ubK4j	  )��}�(h�K2j  ]�h�h�j  K4ubK5j	  )��}�(h�K2j  ]�h�h�j  K5ubK6j	  )��}�(h�K2j  ]�h�h�j  K6ubK7j	  )��}�(h�K2j  ]�h�h�j  K7ubK8j	  )��}�(h�K2j  ]�h�h�j  K8ubK9j	  )��}�(h�K2j  ]�h�h�j  K9ubK:j	  )��}�(h�K2j  ]�h�h�j  K:ubK;j	  )��}�(h�K2j  ]�h�h�j  K;ubK<j	  )��}�(h�K2j  ]�h�h�j  K<ubK=j	  )��}�(h�K2j  ]�h�h�j  K=ubK>j	  )��}�(h�K2j  ]�h�h�j  K>ubK?j	  )��}�(h�K2j  ]�h�h�j  K?ubK@j	  )��}�(h�K2j  ]�h�h�j  K@ubKAj	  )��}�(h�K2j  ]�h�h�j  KAubKBj	  )��}�(h�K2j  ]�h�h�j  KBubKCj	  )��}�(h�K2j  ]�h�h�j  KCubuK3}�(K j	  )��}�(h�K3j  ]�h�h�j  K ubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubK	j	  )��}�(h�K3j  ]�h�h�j  K	ubK
j	  )��}�(h�K3j  ]�h�h�j  K
ubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubKj	  )��}�(h�K3j  ]�h�h�j  KubK j	  )��}�(h�K3j  ]�h�h�j  K ubK!j	  )��}�(h�K3j  ]�h�h�j  K!ubK"j	  )��}�(h�K3j  ]�h�h�j  K"ubK#j	  )��}�(h�K3j  ]�h�h�j  K#ubK$j	  )��}�(h�K3j  ]�h�h�j  K$ubK%j	  )��}�(h�K3j  ]�h�h�j  K%ubK&j	  )��}�(h�K3j  ]�h�h�j  K&ubK'j	  )��}�(h�K3j  ]�h�h�j  K'ubK(j	  )��}�(h�K3j  ]�h�h�j  K(ubK)j	  )��}�(h�K3j  ]�h�h�j  K)ubK*j	  )��}�(h�K3j  ]�h�h�j  K*ubK+j	  )��}�(h�K3j  ]�h�h�j  K+ubK,j	  )��}�(h�K3j  ]�h�h�j  K,ubK-j	  )��}�(h�K3j  ]�h�h�j  K-ubK.j	  )��}�(h�K3j  ]�h�h�j  K.ubK/j	  )��}�(h�K3j  ]�h�h�j  K/ubK0j	  )��}�(h�K3j  ]�h�h�j  K0ubK1j	  )��}�(h�K3j  ]�h�h�j  K1ubK2j	  )��}�(h�K3j  ]�h�h�j  K2ubK3j	  )��}�(h�K3j  ]�h�h�j  K3ubK4j	  )��}�(h�K3j  ]�h�h�j  K4ubK5j	  )��}�(h�K3j  ]�h�h�j  K5ubK6j	  )��}�(h�K3j  ]�h�h�j  K6ubK7j	  )��}�(h�K3j  ]�h�h�j  K7ubK8j	  )��}�(h�K3j  ]�h�h�j  K8ubK9j	  )��}�(h�K3j  ]�h�h�j  K9ubK:j	  )��}�(h�K3j  ]�h�h�j  K:ubK;j	  )��}�(h�K3j  ]�h�h�j  K;ubK<j	  )��}�(h�K3j  ]�h�h�j  K<ubK=j	  )��}�(h�K3j  ]�h�h�j  K=ubK>j	  )��}�(h�K3j  ]�h�h�j  K>ubK?j	  )��}�(h�K3j  ]�h�h�j  K?ubK@j	  )��}�(h�K3j  ]�h�h�j  K@ubKAj	  )��}�(h�K3j  ]�h�h�j  KAubKBj	  )��}�(h�K3j  ]�h�h�j  KBubKCj	  )��}�(h�K3j  ]�h�h�j  KCubuK4}�(K j	  )��}�(h�K4j  ]�h�h�j  K ubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubK	j	  )��}�(h�K4j  ]�h�h�j  K	ubK
j	  )��}�(h�K4j  ]�h�h�j  K
ubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubKj	  )��}�(h�K4j  ]�h�h�j  KubK j	  )��}�(h�K4j  ]�h�h�j  K ubK!j	  )��}�(h�K4j  ]�h�h�j  K!ubK"j	  )��}�(h�K4j  ]�h�h�j  K"ubK#j	  )��}�(h�K4j  ]�h�h�j  K#ubK$j	  )��}�(h�K4j  ]�h�h�j  K$ubK%j	  )��}�(h�K4j  ]�h�h�j  K%ubK&j	  )��}�(h�K4j  ]�h�h�j  K&ubK'j	  )��}�(h�K4j  ]�h�h�j  K'ubK(j	  )��}�(h�K4j  ]�h�h�j  K(ubK)j	  )��}�(h�K4j  ]�h�h�j  K)ubK*j	  )��}�(h�K4j  ]�h�h�j  K*ubK+j	  )��}�(h�K4j  ]�h�h�j  K+ubK,j	  )��}�(h�K4j  ]�h�h�j  K,ubK-j	  )��}�(h�K4j  ]�h�h�j  K-ubK.j	  )��}�(h�K4j  ]�h�h�j  K.ubK/j	  )��}�(h�K4j  ]�h�h�j  K/ubK0j	  )��}�(h�K4j  ]�h�h�j  K0ubK1j	  )��}�(h�K4j  ]�h�h�j  K1ubK2j	  )��}�(h�K4j  ]�h�h�j  K2ubK3j	  )��}�(h�K4j  ]�h�h�j  K3ubK4j	  )��}�(h�K4j  ]�h�h�j  K4ubK5j	  )��}�(h�K4j  ]�h�h�j  K5ubK6j	  )��}�(h�K4j  ]�h�h�j  K6ubK7j	  )��}�(h�K4j  ]�h�h�j  K7ubK8j	  )��}�(h�K4j  ]�h�h�j  K8ubK9j	  )��}�(h�K4j  ]�h�h�j  K9ubK:j	  )��}�(h�K4j  ]�h�h�j  K:ubK;j	  )��}�(h�K4j  ]�h�h�j  K;ubK<j	  )��}�(h�K4j  ]�h�h�j  K<ubK=j	  )��}�(h�K4j  ]�h�h�j  K=ubK>j	  )��}�(h�K4j  ]�h�h�j  K>ubK?j	  )��}�(h�K4j  ]�h�h�j  K?ubK@j	  )��}�(h�K4j  ]�h�h�j  K@ubKAj	  )��}�(h�K4j  ]�h�h�j  KAubKBj	  )��}�(h�K4j  ]�h�h�j  KBubKCj	  )��}�(h�K4j  ]�h�h�j  KCubuK5}�(K j	  )��}�(h�K5j  ]�h�h�j  K ubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubK	j	  )��}�(h�K5j  ]�h�h�j  K	ubK
j	  )��}�(h�K5j  ]�h�h�j  K
ubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubKj	  )��}�(h�K5j  ]�h�h�j  KubK j	  )��}�(h�K5j  ]�h�h�j  K ubK!j	  )��}�(h�K5j  ]�h�h�j  K!ubK"j	  )��}�(h�K5j  ]�h�h�j  K"ubK#j	  )��}�(h�K5j  ]�h�h�j  K#ubK$j	  )��}�(h�K5j  ]�h�h�j  K$ubK%j	  )��}�(h�K5j  ]�h�h�j  K%ubK&j	  )��}�(h�K5j  ]�h�h�j  K&ubK'j	  )��}�(h�K5j  ]�h�h�j  K'ubK(j	  )��}�(h�K5j  ]�h�h�j  K(ubK)j	  )��}�(h�K5j  ]�h�h�j  K)ubK*j	  )��}�(h�K5j  ]�h�h�j  K*ubK+j	  )��}�(h�K5j  ]�h�h�j  K+ubK,j	  )��}�(h�K5j  ]�h�h�j  K,ubK-j	  )��}�(h�K5j  ]�h�h�j  K-ubK.j	  )��}�(h�K5j  ]�h�h�j  K.ubK/j	  )��}�(h�K5j  ]�h�h�j  K/ubK0j	  )��}�(h�K5j  ]�h�h�j  K0ubK1j	  )��}�(h�K5j  ]�h�h�j  K1ubK2j	  )��}�(h�K5j  ]�h�h�j  K2ubK3j	  )��}�(h�K5j  ]�h�h�j  K3ubK4j	  )��}�(h�K5j  ]�h�h�j  K4ubK5j	  )��}�(h�K5j  ]�h�h�j  K5ubK6j	  )��}�(h�K5j  ]�h�h�j  K6ubK7j	  )��}�(h�K5j  ]�h�h�j  K7ubK8j	  )��}�(h�K5j  ]�h�h�j  K8ubK9j	  )��}�(h�K5j  ]�h�h�j  K9ubK:j	  )��}�(h�K5j  ]�h�h�j  K:ubK;j	  )��}�(h�K5j  ]�h�h�j  K;ubK<j	  )��}�(h�K5j  ]�h�h�j  K<ubK=j	  )��}�(h�K5j  ]�Kah�h�j  K=ubK>j	  )��}�(h�K5j  ]�h�h�j  K>ubK?j	  )��}�(h�K5j  ]�h�h�j  K?ubK@j	  )��}�(h�K5j  ]�h�h�j  K@ubKAj	  )��}�(h�K5j  ]�h�h�j  KAubKBj	  )��}�(h�K5j  ]�h�h�j  KBubKCj	  )��}�(h�K5j  ]�h�h�j  KCubuK6}�(K j	  )��}�(h�K6j  ]�h�h�j  K ubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubK	j	  )��}�(h�K6j  ]�h�h�j  K	ubK
j	  )��}�(h�K6j  ]�h�h�j  K
ubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubKj	  )��}�(h�K6j  ]�h�h�j  KubK j	  )��}�(h�K6j  ]�h�h�j  K ubK!j	  )��}�(h�K6j  ]�h�h�j  K!ubK"j	  )��}�(h�K6j  ]�h�h�j  K"ubK#j	  )��}�(h�K6j  ]�h�h�j  K#ubK$j	  )��}�(h�K6j  ]�h�h�j  K$ubK%j	  )��}�(h�K6j  ]�h�h�j  K%ubK&j	  )��}�(h�K6j  ]�h�h�j  K&ubK'j	  )��}�(h�K6j  ]�h�h�j  K'ubK(j	  )��}�(h�K6j  ]�h�h�j  K(ubK)j	  )��}�(h�K6j  ]�h�h�j  K)ubK*j	  )��}�(h�K6j  ]�h�h�j  K*ubK+j	  )��}�(h�K6j  ]�h�h�j  K+ubK,j	  )��}�(h�K6j  ]�h�h�j  K,ubK-j	  )��}�(h�K6j  ]�h�h�j  K-ubK.j	  )��}�(h�K6j  ]�h�h�j  K.ubK/j	  )��}�(h�K6j  ]�h�h�j  K/ubK0j	  )��}�(h�K6j  ]�h�h�j  K0ubK1j	  )��}�(h�K6j  ]�h�h�j  K1ubK2j	  )��}�(h�K6j  ]�h�h�j  K2ubK3j	  )��}�(h�K6j  ]�h�h�j  K3ubK4j	  )��}�(h�K6j  ]�h�h�j  K4ubK5j	  )��}�(h�K6j  ]�h�h�j  K5ubK6j	  )��}�(h�K6j  ]�h�h�j  K6ubK7j	  )��}�(h�K6j  ]�h�h�j  K7ubK8j	  )��}�(h�K6j  ]�h�h�j  K8ubK9j	  )��}�(h�K6j  ]�h�h�j  K9ubK:j	  )��}�(h�K6j  ]�h�h�j  K:ubK;j	  )��}�(h�K6j  ]�h�h�j  K;ubK<j	  )��}�(h�K6j  ]�h�h�j  K<ubK=j	  )��}�(h�K6j  ]�h�h�j  K=ubK>j	  )��}�(h�K6j  ]�h�h�j  K>ubK?j	  )��}�(h�K6j  ]�h�h�j  K?ubK@j	  )��}�(h�K6j  ]�h�h�j  K@ubKAj	  )��}�(h�K6j  ]�h�h�j  KAubKBj	  )��}�(h�K6j  ]�h�h�j  KBubKCj	  )��}�(h�K6j  ]�h�h�j  KCubuK7}�(K j	  )��}�(h�K7j  ]�h�h�j  K ubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubK	j	  )��}�(h�K7j  ]�h�h�j  K	ubK
j	  )��}�(h�K7j  ]�h�h�j  K
ubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubKj	  )��}�(h�K7j  ]�h�h�j  KubK j	  )��}�(h�K7j  ]�h�h�j  K ubK!j	  )��}�(h�K7j  ]�h�h�j  K!ubK"j	  )��}�(h�K7j  ]�h�h�j  K"ubK#j	  )��}�(h�K7j  ]�h�h�j  K#ubK$j	  )��}�(h�K7j  ]�h�h�j  K$ubK%j	  )��}�(h�K7j  ]�h�h�j  K%ubK&j	  )��}�(h�K7j  ]�h�h�j  K&ubK'j	  )��}�(h�K7j  ]�h�h�j  K'ubK(j	  )��}�(h�K7j  ]�h�h�j  K(ubK)j	  )��}�(h�K7j  ]�h�h�j  K)ubK*j	  )��}�(h�K7j  ]�h�h�j  K*ubK+j	  )��}�(h�K7j  ]�h�h�j  K+ubK,j	  )��}�(h�K7j  ]�h�h�j  K,ubK-j	  )��}�(h�K7j  ]�h�h�j  K-ubK.j	  )��}�(h�K7j  ]�h�h�j  K.ubK/j	  )��}�(h�K7j  ]�h�h�j  K/ubK0j	  )��}�(h�K7j  ]�h�h�j  K0ubK1j	  )��}�(h�K7j  ]�h�h�j  K1ubK2j	  )��}�(h�K7j  ]�h�h�j  K2ubK3j	  )��}�(h�K7j  ]�h�h�j  K3ubK4j	  )��}�(h�K7j  ]�h�h�j  K4ubK5j	  )��}�(h�K7j  ]�h�h�j  K5ubK6j	  )��}�(h�K7j  ]�h�h�j  K6ubK7j	  )��}�(h�K7j  ]�h�h�j  K7ubK8j	  )��}�(h�K7j  ]�h�h�j  K8ubK9j	  )��}�(h�K7j  ]�h�h�j  K9ubK:j	  )��}�(h�K7j  ]�h�h�j  K:ubK;j	  )��}�(h�K7j  ]�h�h�j  K;ubK<j	  )��}�(h�K7j  ]�h�h�j  K<ubK=j	  )��}�(h�K7j  ]�Kah�h�j  K=ubK>j	  )��}�(h�K7j  ]�h�h�j  K>ubK?j	  )��}�(h�K7j  ]�h�h�j  K?ubK@j	  )��}�(h�K7j  ]�Kah�h�j  K@ubKAj	  )��}�(h�K7j  ]�h�h�j  KAubKBj	  )��}�(h�K7j  ]�h�h�j  KBubKCj	  )��}�(h�K7j  ]�h�h�j  KCubuK8}�(K j	  )��}�(h�K8j  ]�h�h�j  K ubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubK	j	  )��}�(h�K8j  ]�h�h�j  K	ubK
j	  )��}�(h�K8j  ]�h�h�j  K
ubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubKj	  )��}�(h�K8j  ]�h�h�j  KubK j	  )��}�(h�K8j  ]�h�h�j  K ubK!j	  )��}�(h�K8j  ]�h�h�j  K!ubK"j	  )��}�(h�K8j  ]�h�h�j  K"ubK#j	  )��}�(h�K8j  ]�h�h�j  K#ubK$j	  )��}�(h�K8j  ]�h�h�j  K$ubK%j	  )��}�(h�K8j  ]�h�h�j  K%ubK&j	  )��}�(h�K8j  ]�h�h�j  K&ubK'j	  )��}�(h�K8j  ]�h�h�j  K'ubK(j	  )��}�(h�K8j  ]�h�h�j  K(ubK)j	  )��}�(h�K8j  ]�h�h�j  K)ubK*j	  )��}�(h�K8j  ]�h�h�j  K*ubK+j	  )��}�(h�K8j  ]�h�h�j  K+ubK,j	  )��}�(h�K8j  ]�h�h�j  K,ubK-j	  )��}�(h�K8j  ]�h�h�j  K-ubK.j	  )��}�(h�K8j  ]�h�h�j  K.ubK/j	  )��}�(h�K8j  ]�h�h�j  K/ubK0j	  )��}�(h�K8j  ]�h�h�j  K0ubK1j	  )��}�(h�K8j  ]�h�h�j  K1ubK2j	  )��}�(h�K8j  ]�h�h�j  K2ubK3j	  )��}�(h�K8j  ]�h�h�j  K3ubK4j	  )��}�(h�K8j  ]�h�h�j  K4ubK5j	  )��}�(h�K8j  ]�h�h�j  K5ubK6j	  )��}�(h�K8j  ]�h�h�j  K6ubK7j	  )��}�(h�K8j  ]�h�h�j  K7ubK8j	  )��}�(h�K8j  ]�h�h�j  K8ubK9j	  )��}�(h�K8j  ]�h�h�j  K9ubK:j	  )��}�(h�K8j  ]�h�h�j  K:ubK;j	  )��}�(h�K8j  ]�h�h�j  K;ubK<j	  )��}�(h�K8j  ]�h�h�j  K<ubK=j	  )��}�(h�K8j  ]�h�h�j  K=ubK>j	  )��}�(h�K8j  ]�h�h�j  K>ubK?j	  )��}�(h�K8j  ]�h�h�j  K?ubK@j	  )��}�(h�K8j  ]�h�h�j  K@ubKAj	  )��}�(h�K8j  ]�h�h�j  KAubKBj	  )��}�(h�K8j  ]�h�h�j  KBubKCj	  )��}�(h�K8j  ]�h�h�j  KCubuK9}�(K j	  )��}�(h�K9j  ]�h�h�j  K ubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubK	j	  )��}�(h�K9j  ]�h�h�j  K	ubK
j	  )��}�(h�K9j  ]�h�h�j  K
ubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubKj	  )��}�(h�K9j  ]�h�h�j  KubK j	  )��}�(h�K9j  ]�h�h�j  K ubK!j	  )��}�(h�K9j  ]�h�h�j  K!ubK"j	  )��}�(h�K9j  ]�h�h�j  K"ubK#j	  )��}�(h�K9j  ]�h�h�j  K#ubK$j	  )��}�(h�K9j  ]�h�h�j  K$ubK%j	  )��}�(h�K9j  ]�h�h�j  K%ubK&j	  )��}�(h�K9j  ]�h�h�j  K&ubK'j	  )��}�(h�K9j  ]�h�h�j  K'ubK(j	  )��}�(h�K9j  ]�h�h�j  K(ubK)j	  )��}�(h�K9j  ]�h�h�j  K)ubK*j	  )��}�(h�K9j  ]�h�h�j  K*ubK+j	  )��}�(h�K9j  ]�h�h�j  K+ubK,j	  )��}�(h�K9j  ]�h�h�j  K,ubK-j	  )��}�(h�K9j  ]�h�h�j  K-ubK.j	  )��}�(h�K9j  ]�h�h�j  K.ubK/j	  )��}�(h�K9j  ]�h�h�j  K/ubK0j	  )��}�(h�K9j  ]�h�h�j  K0ubK1j	  )��}�(h�K9j  ]�h�h�j  K1ubK2j	  )��}�(h�K9j  ]�h�h�j  K2ubK3j	  )��}�(h�K9j  ]�h�h�j  K3ubK4j	  )��}�(h�K9j  ]�h�h�j  K4ubK5j	  )��}�(h�K9j  ]�h�h�j  K5ubK6j	  )��}�(h�K9j  ]�h�h�j  K6ubK7j	  )��}�(h�K9j  ]�h�h�j  K7ubK8j	  )��}�(h�K9j  ]�h�h�j  K8ubK9j	  )��}�(h�K9j  ]�h�h�j  K9ubK:j	  )��}�(h�K9j  ]�h�h�j  K:ubK;j	  )��}�(h�K9j  ]�h�h�j  K;ubK<j	  )��}�(h�K9j  ]�h�h�j  K<ubK=j	  )��}�(h�K9j  ]�h�h�j  K=ubK>j	  )��}�(h�K9j  ]�h�h�j  K>ubK?j	  )��}�(h�K9j  ]�h�h�j  K?ubK@j	  )��}�(h�K9j  ]�h�h�j  K@ubKAj	  )��}�(h�K9j  ]�h�h�j  KAubKBj	  )��}�(h�K9j  ]�h�h�j  KBubKCj	  )��}�(h�K9j  ]�h�h�j  KCubuK:}�(K j	  )��}�(h�K:j  ]�h�h�j  K ubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubK	j	  )��}�(h�K:j  ]�h�h�j  K	ubK
j	  )��}�(h�K:j  ]�h�h�j  K
ubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubKj	  )��}�(h�K:j  ]�h�h�j  KubK j	  )��}�(h�K:j  ]�h�h�j  K ubK!j	  )��}�(h�K:j  ]�h�h�j  K!ubK"j	  )��}�(h�K:j  ]�h�h�j  K"ubK#j	  )��}�(h�K:j  ]�h�h�j  K#ubK$j	  )��}�(h�K:j  ]�h�h�j  K$ubK%j	  )��}�(h�K:j  ]�h�h�j  K%ubK&j	  )��}�(h�K:j  ]�h�h�j  K&ubK'j	  )��}�(h�K:j  ]�h�h�j  K'ubK(j	  )��}�(h�K:j  ]�h�h�j  K(ubK)j	  )��}�(h�K:j  ]�h�h�j  K)ubK*j	  )��}�(h�K:j  ]�h�h�j  K*ubK+j	  )��}�(h�K:j  ]�h�h�j  K+ubK,j	  )��}�(h�K:j  ]�h�h�j  K,ubK-j	  )��}�(h�K:j  ]�h�h�j  K-ubK.j	  )��}�(h�K:j  ]�h�h�j  K.ubK/j	  )��}�(h�K:j  ]�h�h�j  K/ubK0j	  )��}�(h�K:j  ]�h�h�j  K0ubK1j	  )��}�(h�K:j  ]�h�h�j  K1ubK2j	  )��}�(h�K:j  ]�h�h�j  K2ubK3j	  )��}�(h�K:j  ]�h�h�j  K3ubK4j	  )��}�(h�K:j  ]�h�h�j  K4ubK5j	  )��}�(h�K:j  ]�h�h�j  K5ubK6j	  )��}�(h�K:j  ]�h�h�j  K6ubK7j	  )��}�(h�K:j  ]�h�h�j  K7ubK8j	  )��}�(h�K:j  ]�h�h�j  K8ubK9j	  )��}�(h�K:j  ]�h�h�j  K9ubK:j	  )��}�(h�K:j  ]�h�h�j  K:ubK;j	  )��}�(h�K:j  ]�h�h�j  K;ubK<j	  )��}�(h�K:j  ]�h�h�j  K<ubK=j	  )��}�(h�K:j  ]�h�h�j  K=ubK>j	  )��}�(h�K:j  ]�h�h�j  K>ubK?j	  )��}�(h�K:j  ]�h�h�j  K?ubK@j	  )��}�(h�K:j  ]�h�h�j  K@ubKAj	  )��}�(h�K:j  ]�h�h�j  KAubKBj	  )��}�(h�K:j  ]�h�h�j  KBubKCj	  )��}�(h�K:j  ]�h�h�j  KCubuK;}�(K j	  )��}�(h�K;j  ]�h�h�j  K ubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�Kah�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubK	j	  )��}�(h�K;j  ]�h�h�j  K	ubK
j	  )��}�(h�K;j  ]�h�h�j  K
ubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubKj	  )��}�(h�K;j  ]�h�h�j  KubK j	  )��}�(h�K;j  ]�h�h�j  K ubK!j	  )��}�(h�K;j  ]�h�h�j  K!ubK"j	  )��}�(h�K;j  ]�h�h�j  K"ubK#j	  )��}�(h�K;j  ]�h�h�j  K#ubK$j	  )��}�(h�K;j  ]�h�h�j  K$ubK%j	  )��}�(h�K;j  ]�h�h�j  K%ubK&j	  )��}�(h�K;j  ]�h�h�j  K&ubK'j	  )��}�(h�K;j  ]�h�h�j  K'ubK(j	  )��}�(h�K;j  ]�h�h�j  K(ubK)j	  )��}�(h�K;j  ]�h�h�j  K)ubK*j	  )��}�(h�K;j  ]�h�h�j  K*ubK+j	  )��}�(h�K;j  ]�h�h�j  K+ubK,j	  )��}�(h�K;j  ]�h�h�j  K,ubK-j	  )��}�(h�K;j  ]�h�h�j  K-ubK.j	  )��}�(h�K;j  ]�h�h�j  K.ubK/j	  )��}�(h�K;j  ]�h�h�j  K/ubK0j	  )��}�(h�K;j  ]�h�h�j  K0ubK1j	  )��}�(h�K;j  ]�h�h�j  K1ubK2j	  )��}�(h�K;j  ]�h�h�j  K2ubK3j	  )��}�(h�K;j  ]�h�h�j  K3ubK4j	  )��}�(h�K;j  ]�h�h�j  K4ubK5j	  )��}�(h�K;j  ]�h�h�j  K5ubK6j	  )��}�(h�K;j  ]�h�h�j  K6ubK7j	  )��}�(h�K;j  ]�h�h�j  K7ubK8j	  )��}�(h�K;j  ]�h�h�j  K8ubK9j	  )��}�(h�K;j  ]�h�h�j  K9ubK:j	  )��}�(h�K;j  ]�h�h�j  K:ubK;j	  )��}�(h�K;j  ]�h�h�j  K;ubK<j	  )��}�(h�K;j  ]�h�h�j  K<ubK=j	  )��}�(h�K;j  ]�h�h�j  K=ubK>j	  )��}�(h�K;j  ]�h�h�j  K>ubK?j	  )��}�(h�K;j  ]�h�h�j  K?ubK@j	  )��}�(h�K;j  ]�h�h�j  K@ubKAj	  )��}�(h�K;j  ]�h�h�j  KAubKBj	  )��}�(h�K;j  ]�h�h�j  KBubKCj	  )��}�(h�K;j  ]�h�h�j  KCubuK<}�(K j	  )��}�(h�K<j  ]�h�h�j  K ubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubK	j	  )��}�(h�K<j  ]�h�h�j  K	ubK
j	  )��}�(h�K<j  ]�h�h�j  K
ubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�Kah�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubKj	  )��}�(h�K<j  ]�h�h�j  KubK j	  )��}�(h�K<j  ]�h�h�j  K ubK!j	  )��}�(h�K<j  ]�h�h�j  K!ubK"j	  )��}�(h�K<j  ]�h�h�j  K"ubK#j	  )��}�(h�K<j  ]�h�h�j  K#ubK$j	  )��}�(h�K<j  ]�h�h�j  K$ubK%j	  )��}�(h�K<j  ]�h�h�j  K%ubK&j	  )��}�(h�K<j  ]�h�h�j  K&ubK'j	  )��}�(h�K<j  ]�h�h�j  K'ubK(j	  )��}�(h�K<j  ]�h�h�j  K(ubK)j	  )��}�(h�K<j  ]�h�h�j  K)ubK*j	  )��}�(h�K<j  ]�h�h�j  K*ubK+j	  )��}�(h�K<j  ]�h�h�j  K+ubK,j	  )��}�(h�K<j  ]�h�h�j  K,ubK-j	  )��}�(h�K<j  ]�h�h�j  K-ubK.j	  )��}�(h�K<j  ]�h�h�j  K.ubK/j	  )��}�(h�K<j  ]�h�h�j  K/ubK0j	  )��}�(h�K<j  ]�h�h�j  K0ubK1j	  )��}�(h�K<j  ]�h�h�j  K1ubK2j	  )��}�(h�K<j  ]�h�h�j  K2ubK3j	  )��}�(h�K<j  ]�h�h�j  K3ubK4j	  )��}�(h�K<j  ]�h�h�j  K4ubK5j	  )��}�(h�K<j  ]�h�h�j  K5ubK6j	  )��}�(h�K<j  ]�h�h�j  K6ubK7j	  )��}�(h�K<j  ]�h�h�j  K7ubK8j	  )��}�(h�K<j  ]�h�h�j  K8ubK9j	  )��}�(h�K<j  ]�h�h�j  K9ubK:j	  )��}�(h�K<j  ]�h�h�j  K:ubK;j	  )��}�(h�K<j  ]�h�h�j  K;ubK<j	  )��}�(h�K<j  ]�h�h�j  K<ubK=j	  )��}�(h�K<j  ]�h�h�j  K=ubK>j	  )��}�(h�K<j  ]�h�h�j  K>ubK?j	  )��}�(h�K<j  ]�h�h�j  K?ubK@j	  )��}�(h�K<j  ]�h�h�j  K@ubKAj	  )��}�(h�K<j  ]�h�h�j  KAubKBj	  )��}�(h�K<j  ]�h�h�j  KBubKCj	  )��}�(h�K<j  ]�h�h�j  KCubuK=}�(K j	  )��}�(h�K=j  ]�h�h�j  K ubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�Kah�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubK	j	  )��}�(h�K=j  ]�h�h�j  K	ubK
j	  )��}�(h�K=j  ]�h�h�j  K
ubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�Kah�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�Kah�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubKj	  )��}�(h�K=j  ]�h�h�j  KubK j	  )��}�(h�K=j  ]�h�h�j  K ubK!j	  )��}�(h�K=j  ]�h�h�j  K!ubK"j	  )��}�(h�K=j  ]�h�h�j  K"ubK#j	  )��}�(h�K=j  ]�h�h�j  K#ubK$j	  )��}�(h�K=j  ]�h�h�j  K$ubK%j	  )��}�(h�K=j  ]�h�h�j  K%ubK&j	  )��}�(h�K=j  ]�h�h�j  K&ubK'j	  )��}�(h�K=j  ]�h�h�j  K'ubK(j	  )��}�(h�K=j  ]�h�h�j  K(ubK)j	  )��}�(h�K=j  ]�h�h�j  K)ubK*j	  )��}�(h�K=j  ]�h�h�j  K*ubK+j	  )��}�(h�K=j  ]�h�h�j  K+ubK,j	  )��}�(h�K=j  ]�h�h�j  K,ubK-j	  )��}�(h�K=j  ]�h�h�j  K-ubK.j	  )��}�(h�K=j  ]�h�h�j  K.ubK/j	  )��}�(h�K=j  ]�h�h�j  K/ubK0j	  )��}�(h�K=j  ]�h�h�j  K0ubK1j	  )��}�(h�K=j  ]�h�h�j  K1ubK2j	  )��}�(h�K=j  ]�h�h�j  K2ubK3j	  )��}�(h�K=j  ]�h�h�j  K3ubK4j	  )��}�(h�K=j  ]�h�h�j  K4ubK5j	  )��}�(h�K=j  ]�h�h�j  K5ubK6j	  )��}�(h�K=j  ]�h�h�j  K6ubK7j	  )��}�(h�K=j  ]�h�h�j  K7ubK8j	  )��}�(h�K=j  ]�h�h�j  K8ubK9j	  )��}�(h�K=j  ]�h�h�j  K9ubK:j	  )��}�(h�K=j  ]�h�h�j  K:ubK;j	  )��}�(h�K=j  ]�h�h�j  K;ubK<j	  )��}�(h�K=j  ]�h�h�j  K<ubK=j	  )��}�(h�K=j  ]�h�h�j  K=ubK>j	  )��}�(h�K=j  ]�h�h�j  K>ubK?j	  )��}�(h�K=j  ]�h�h�j  K?ubK@j	  )��}�(h�K=j  ]�h�h�j  K@ubKAj	  )��}�(h�K=j  ]�h�h�j  KAubKBj	  )��}�(h�K=j  ]�h�h�j  KBubKCj	  )��}�(h�K=j  ]�h�h�j  KCubuK>}�(K j	  )��}�(h�K>j  ]�h�h�j  K ubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�Kah�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubK	j	  )��}�(h�K>j  ]�h�h�j  K	ubK
j	  )��}�(h�K>j  ]�h�h�j  K
ubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�Kah�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubKj	  )��}�(h�K>j  ]�h�h�j  KubK j	  )��}�(h�K>j  ]�h�h�j  K ubK!j	  )��}�(h�K>j  ]�h�h�j  K!ubK"j	  )��}�(h�K>j  ]�h�h�j  K"ubK#j	  )��}�(h�K>j  ]�h�h�j  K#ubK$j	  )��}�(h�K>j  ]�h�h�j  K$ubK%j	  )��}�(h�K>j  ]�h�h�j  K%ubK&j	  )��}�(h�K>j  ]�h�h�j  K&ubK'j	  )��}�(h�K>j  ]�h�h�j  K'ubK(j	  )��}�(h�K>j  ]�h�h�j  K(ubK)j	  )��}�(h�K>j  ]�h�h�j  K)ubK*j	  )��}�(h�K>j  ]�h�h�j  K*ubK+j	  )��}�(h�K>j  ]�h�h�j  K+ubK,j	  )��}�(h�K>j  ]�h�h�j  K,ubK-j	  )��}�(h�K>j  ]�h�h�j  K-ubK.j	  )��}�(h�K>j  ]�h�h�j  K.ubK/j	  )��}�(h�K>j  ]�h�h�j  K/ubK0j	  )��}�(h�K>j  ]�h�h�j  K0ubK1j	  )��}�(h�K>j  ]�h�h�j  K1ubK2j	  )��}�(h�K>j  ]�h�h�j  K2ubK3j	  )��}�(h�K>j  ]�h�h�j  K3ubK4j	  )��}�(h�K>j  ]�h�h�j  K4ubK5j	  )��}�(h�K>j  ]�h�h�j  K5ubK6j	  )��}�(h�K>j  ]�h�h�j  K6ubK7j	  )��}�(h�K>j  ]�h�h�j  K7ubK8j	  )��}�(h�K>j  ]�h�h�j  K8ubK9j	  )��}�(h�K>j  ]�h�h�j  K9ubK:j	  )��}�(h�K>j  ]�h�h�j  K:ubK;j	  )��}�(h�K>j  ]�h�h�j  K;ubK<j	  )��}�(h�K>j  ]�h�h�j  K<ubK=j	  )��}�(h�K>j  ]�h�h�j  K=ubK>j	  )��}�(h�K>j  ]�h�h�j  K>ubK?j	  )��}�(h�K>j  ]�h�h�j  K?ubK@j	  )��}�(h�K>j  ]�h�h�j  K@ubKAj	  )��}�(h�K>j  ]�h�h�j  KAubKBj	  )��}�(h�K>j  ]�h�h�j  KBubKCj	  )��}�(h�K>j  ]�h�h�j  KCubuK?}�(K j	  )��}�(h�K?j  ]�h�h�j  K ubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubK	j	  )��}�(h�K?j  ]�h�h�j  K	ubK
j	  )��}�(h�K?j  ]�h�h�j  K
ubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�Kah�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubKj	  )��}�(h�K?j  ]�h�h�j  KubK j	  )��}�(h�K?j  ]�h�h�j  K ubK!j	  )��}�(h�K?j  ]�h�h�j  K!ubK"j	  )��}�(h�K?j  ]�h�h�j  K"ubK#j	  )��}�(h�K?j  ]�h�h�j  K#ubK$j	  )��}�(h�K?j  ]�h�h�j  K$ubK%j	  )��}�(h�K?j  ]�h�h�j  K%ubK&j	  )��}�(h�K?j  ]�h�h�j  K&ubK'j	  )��}�(h�K?j  ]�Kah�h�j  K'ubK(j	  )��}�(h�K?j  ]�h�h�j  K(ubK)j	  )��}�(h�K?j  ]�h�h�j  K)ubK*j	  )��}�(h�K?j  ]�h�h�j  K*ubK+j	  )��}�(h�K?j  ]�h�h�j  K+ubK,j	  )��}�(h�K?j  ]�h�h�j  K,ubK-j	  )��}�(h�K?j  ]�h�h�j  K-ubK.j	  )��}�(h�K?j  ]�h�h�j  K.ubK/j	  )��}�(h�K?j  ]�h�h�j  K/ubK0j	  )��}�(h�K?j  ]�h�h�j  K0ubK1j	  )��}�(h�K?j  ]�h�h�j  K1ubK2j	  )��}�(h�K?j  ]�h�h�j  K2ubK3j	  )��}�(h�K?j  ]�h�h�j  K3ubK4j	  )��}�(h�K?j  ]�h�h�j  K4ubK5j	  )��}�(h�K?j  ]�h�h�j  K5ubK6j	  )��}�(h�K?j  ]�h�h�j  K6ubK7j	  )��}�(h�K?j  ]�h�h�j  K7ubK8j	  )��}�(h�K?j  ]�h�h�j  K8ubK9j	  )��}�(h�K?j  ]�h�h�j  K9ubK:j	  )��}�(h�K?j  ]�h�h�j  K:ubK;j	  )��}�(h�K?j  ]�h�h�j  K;ubK<j	  )��}�(h�K?j  ]�h�h�j  K<ubK=j	  )��}�(h�K?j  ]�h�h�j  K=ubK>j	  )��}�(h�K?j  ]�h�h�j  K>ubK?j	  )��}�(h�K?j  ]�h�h�j  K?ubK@j	  )��}�(h�K?j  ]�h�h�j  K@ubKAj	  )��}�(h�K?j  ]�h�h�j  KAubKBj	  )��}�(h�K?j  ]�h�h�j  KBubKCj	  )��}�(h�K?j  ]�h�h�j  KCubuK@}�(K j	  )��}�(h�K@j  ]�h�h�j  K ubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubK	j	  )��}�(h�K@j  ]�h�h�j  K	ubK
j	  )��}�(h�K@j  ]�h�h�j  K
ubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubKj	  )��}�(h�K@j  ]�h�h�j  KubK j	  )��}�(h�K@j  ]�h�h�j  K ubK!j	  )��}�(h�K@j  ]�h�h�j  K!ubK"j	  )��}�(h�K@j  ]�h�h�j  K"ubK#j	  )��}�(h�K@j  ]�h�h�j  K#ubK$j	  )��}�(h�K@j  ]�Kah�h�j  K$ubK%j	  )��}�(h�K@j  ]�Kah�h�j  K%ubK&j	  )��}�(h�K@j  ]�h�h�j  K&ubK'j	  )��}�(h�K@j  ]�h�h�j  K'ubK(j	  )��}�(h�K@j  ]�h�h�j  K(ubK)j	  )��}�(h�K@j  ]�h�h�j  K)ubK*j	  )��}�(h�K@j  ]�h�h�j  K*ubK+j	  )��}�(h�K@j  ]�h�h�j  K+ubK,j	  )��}�(h�K@j  ]�h�h�j  K,ubK-j	  )��}�(h�K@j  ]�h�h�j  K-ubK.j	  )��}�(h�K@j  ]�h�h�j  K.ubK/j	  )��}�(h�K@j  ]�h�h�j  K/ubK0j	  )��}�(h�K@j  ]�h�h�j  K0ubK1j	  )��}�(h�K@j  ]�h�h�j  K1ubK2j	  )��}�(h�K@j  ]�h�h�j  K2ubK3j	  )��}�(h�K@j  ]�h�h�j  K3ubK4j	  )��}�(h�K@j  ]�h�h�j  K4ubK5j	  )��}�(h�K@j  ]�h�h�j  K5ubK6j	  )��}�(h�K@j  ]�h�h�j  K6ubK7j	  )��}�(h�K@j  ]�h�h�j  K7ubK8j	  )��}�(h�K@j  ]�h�h�j  K8ubK9j	  )��}�(h�K@j  ]�h�h�j  K9ubK:j	  )��}�(h�K@j  ]�h�h�j  K:ubK;j	  )��}�(h�K@j  ]�h�h�j  K;ubK<j	  )��}�(h�K@j  ]�h�h�j  K<ubK=j	  )��}�(h�K@j  ]�h�h�j  K=ubK>j	  )��}�(h�K@j  ]�h�h�j  K>ubK?j	  )��}�(h�K@j  ]�h�h�j  K?ubK@j	  )��}�(h�K@j  ]�h�h�j  K@ubKAj	  )��}�(h�K@j  ]�h�h�j  KAubKBj	  )��}�(h�K@j  ]�h�h�j  KBubKCj	  )��}�(h�K@j  ]�h�h�j  KCubuKA}�(K j	  )��}�(h�KAj  ]�h�h�j  K ubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubK	j	  )��}�(h�KAj  ]�h�h�j  K	ubK
j	  )��}�(h�KAj  ]�h�h�j  K
ubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubKj	  )��}�(h�KAj  ]�h�h�j  KubK j	  )��}�(h�KAj  ]�h�h�j  K ubK!j	  )��}�(h�KAj  ]�h�h�j  K!ubK"j	  )��}�(h�KAj  ]�Kah�h�j  K"ubK#j	  )��}�(h�KAj  ]�h�h�j  K#ubK$j	  )��}�(h�KAj  ]�h�h�j  K$ubK%j	  )��}�(h�KAj  ]�h�h�j  K%ubK&j	  )��}�(h�KAj  ]�h�h�j  K&ubK'j	  )��}�(h�KAj  ]�h�h�j  K'ubK(j	  )��}�(h�KAj  ]�h�h�j  K(ubK)j	  )��}�(h�KAj  ]�h�h�j  K)ubK*j	  )��}�(h�KAj  ]�h�h�j  K*ubK+j	  )��}�(h�KAj  ]�h�h�j  K+ubK,j	  )��}�(h�KAj  ]�h�h�j  K,ubK-j	  )��}�(h�KAj  ]�h�h�j  K-ubK.j	  )��}�(h�KAj  ]�h�h�j  K.ubK/j	  )��}�(h�KAj  ]�h�h�j  K/ubK0j	  )��}�(h�KAj  ]�h�h�j  K0ubK1j	  )��}�(h�KAj  ]�h�h�j  K1ubK2j	  )��}�(h�KAj  ]�h�h�j  K2ubK3j	  )��}�(h�KAj  ]�h�h�j  K3ubK4j	  )��}�(h�KAj  ]�h�h�j  K4ubK5j	  )��}�(h�KAj  ]�h�h�j  K5ubK6j	  )��}�(h�KAj  ]�h�h�j  K6ubK7j	  )��}�(h�KAj  ]�h�h�j  K7ubK8j	  )��}�(h�KAj  ]�h�h�j  K8ubK9j	  )��}�(h�KAj  ]�h�h�j  K9ubK:j	  )��}�(h�KAj  ]�h�h�j  K:ubK;j	  )��}�(h�KAj  ]�h�h�j  K;ubK<j	  )��}�(h�KAj  ]�h�h�j  K<ubK=j	  )��}�(h�KAj  ]�h�h�j  K=ubK>j	  )��}�(h�KAj  ]�h�h�j  K>ubK?j	  )��}�(h�KAj  ]�h�h�j  K?ubK@j	  )��}�(h�KAj  ]�h�h�j  K@ubKAj	  )��}�(h�KAj  ]�h�h�j  KAubKBj	  )��}�(h�KAj  ]�h�h�j  KBubKCj	  )��}�(h�KAj  ]�h�h�j  KCubuKB}�(K j	  )��}�(h�KBj  ]�h�h�j  K ubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubK	j	  )��}�(h�KBj  ]�h�h�j  K	ubK
j	  )��}�(h�KBj  ]�h�h�j  K
ubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubKj	  )��}�(h�KBj  ]�h�h�j  KubK j	  )��}�(h�KBj  ]�h�h�j  K ubK!j	  )��}�(h�KBj  ]�h�h�j  K!ubK"j	  )��}�(h�KBj  ]�h�h�j  K"ubK#j	  )��}�(h�KBj  ]�h�h�j  K#ubK$j	  )��}�(h�KBj  ]�h�h�j  K$ubK%j	  )��}�(h�KBj  ]�h�h�j  K%ubK&j	  )��}�(h�KBj  ]�h�h�j  K&ubK'j	  )��}�(h�KBj  ]�h�h�j  K'ubK(j	  )��}�(h�KBj  ]�h�h�j  K(ubK)j	  )��}�(h�KBj  ]�h�h�j  K)ubK*j	  )��}�(h�KBj  ]�h�h�j  K*ubK+j	  )��}�(h�KBj  ]�h�h�j  K+ubK,j	  )��}�(h�KBj  ]�h�h�j  K,ubK-j	  )��}�(h�KBj  ]�h�h�j  K-ubK.j	  )��}�(h�KBj  ]�h�h�j  K.ubK/j	  )��}�(h�KBj  ]�h�h�j  K/ubK0j	  )��}�(h�KBj  ]�h�h�j  K0ubK1j	  )��}�(h�KBj  ]�h�h�j  K1ubK2j	  )��}�(h�KBj  ]�h�h�j  K2ubK3j	  )��}�(h�KBj  ]�h�h�j  K3ubK4j	  )��}�(h�KBj  ]�h�h�j  K4ubK5j	  )��}�(h�KBj  ]�h�h�j  K5ubK6j	  )��}�(h�KBj  ]�h�h�j  K6ubK7j	  )��}�(h�KBj  ]�h�h�j  K7ubK8j	  )��}�(h�KBj  ]�h�h�j  K8ubK9j	  )��}�(h�KBj  ]�h�h�j  K9ubK:j	  )��}�(h�KBj  ]�h�h�j  K:ubK;j	  )��}�(h�KBj  ]�h�h�j  K;ubK<j	  )��}�(h�KBj  ]�h�h�j  K<ubK=j	  )��}�(h�KBj  ]�h�h�j  K=ubK>j	  )��}�(h�KBj  ]�h�h�j  K>ubK?j	  )��}�(h�KBj  ]�h�h�j  K?ubK@j	  )��}�(h�KBj  ]�h�h�j  K@ubKAj	  )��}�(h�KBj  ]�h�h�j  KAubKBj	  )��}�(h�KBj  ]�h�h�j  KBubKCj	  )��}�(h�KBj  ]�h�h�j  KCubuKC}�(K j	  )��}�(h�KCj  ]�h�h�j  K ubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubK	j	  )��}�(h�KCj  ]�h�h�j  K	ubK
j	  )��}�(h�KCj  ]�h�h�j  K
ubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubKj	  )��}�(h�KCj  ]�h�h�j  KubK j	  )��}�(h�KCj  ]�h�h�j  K ubK!j	  )��}�(h�KCj  ]�h�h�j  K!ubK"j	  )��}�(h�KCj  ]�h�h�j  K"ubK#j	  )��}�(h�KCj  ]�h�h�j  K#ubK$j	  )��}�(h�KCj  ]�h�h�j  K$ubK%j	  )��}�(h�KCj  ]�h�h�j  K%ubK&j	  )��}�(h�KCj  ]�h�h�j  K&ubK'j	  )��}�(h�KCj  ]�h�h�j  K'ubK(j	  )��}�(h�KCj  ]�h�h�j  K(ubK)j	  )��}�(h�KCj  ]�h�h�j  K)ubK*j	  )��}�(h�KCj  ]�h�h�j  K*ubK+j	  )��}�(h�KCj  ]�h�h�j  K+ubK,j	  )��}�(h�KCj  ]�h�h�j  K,ubK-j	  )��}�(h�KCj  ]�h�h�j  K-ubK.j	  )��}�(h�KCj  ]�h�h�j  K.ubK/j	  )��}�(h�KCj  ]�h�h�j  K/ubK0j	  )��}�(h�KCj  ]�h�h�j  K0ubK1j	  )��}�(h�KCj  ]�h�h�j  K1ubK2j	  )��}�(h�KCj  ]�h�h�j  K2ubK3j	  )��}�(h�KCj  ]�h�h�j  K3ubK4j	  )��}�(h�KCj  ]�h�h�j  K4ubK5j	  )��}�(h�KCj  ]�h�h�j  K5ubK6j	  )��}�(h�KCj  ]�h�h�j  K6ubK7j	  )��}�(h�KCj  ]�h�h�j  K7ubK8j	  )��}�(h�KCj  ]�h�h�j  K8ubK9j	  )��}�(h�KCj  ]�h�h�j  K9ubK:j	  )��}�(h�KCj  ]�h�h�j  K:ubK;j	  )��}�(h�KCj  ]�h�h�j  K;ubK<j	  )��}�(h�KCj  ]�h�h�j  K<ubK=j	  )��}�(h�KCj  ]�h�h�j  K=ubK>j	  )��}�(h�KCj  ]�h�h�j  K>ubK?j	  )��}�(h�KCj  ]�h�h�j  K?ubK@j	  )��}�(h�KCj  ]�h�h�j  K@ubKAj	  )��}�(h�KCj  ]�h�h�j  KAubKBj	  )��}�(h�KCj  ]�h�h�j  KBubKCj	  )��}�(h�KCj  ]�h�h�j  KCubuu�	tilesSeen�]��djikstra_Stairs_Down�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NKaK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKGKFKEKFKEKDKEKFKGKHKIKJKKKLKMKNKOKPKQKRKSKTKSKTKUKVKWKXKYKZK[K\K]K^K_K`KaKbNe]�(NK`K_K^K]NNKZKYKXKWKVKUKTKSKRKQKPKOKNNKLKKKJKIKHKGKFKEKFKEKDKEKDKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQKRKSKRKSKTKUKVKWKXNKZK[K\K]K^NK`KaNe]�(NK_K^K]K\K[NKYKXKWKVKUNNKRNKPKOKNKMKLKKNKIKHKGKFKEKDKEKDKCKDKCKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQKRKQKRKSKTKUKVKWKXKYKZK[K\K]K^K_K`Ne]�(NK^K]K\NKZKYKXKWNKUKTKSKRKQNKOKNKMKLKKKJKIKHKGKFKEKDKCKDKCKBKCKBKAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQKPKQKRKSKTKUKVKWKXKYKZK[K\K]K^K_Ne]�(NK]K\K[NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKCKBKAKBKAK@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKONKOKPNKTKSKTKUKVKWKXKYNK[K\K]K^Ne]�(NK\K[KZKYKXKWKVKUKTKSKRKQKPNKNKMKLKKKJKIKHKGKFKEKDKCKBKAKBKAK@KAK@K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNNKNKOKPNKRKSKTKUKVKWKXKYKZNK\K]Ne]�(NK[KZKYKXKWKVKUKTKSKRNKPKOKNKMKLKKNKINKGKFKEKDKCKBKAK@KAK@K?K@K?K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMNKMKNKOKPKQKRKSKTKUKVKWKXKYKZK[K\Ne]�(NKZKYNKWKVKUKTKSKRKQKPKONKMKLNKJKIKHKGKFKEKDKCKBKAK@K?K@K?K>K?K>K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKKKLKMNKOKPNKRKSKTKUKVKWKXKYKZK[Ne]�(NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKHNKDKCNNK@K?K>K?K>K=K>K=K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKJKKKLKMKNKONKQKRKSKTKUKVNKXKYKZNe]�(NKXKWKVKUKTKUKTNKPKOKNKMKLNKJKIKHKGKFNKDNKBKAK@K?K>K=NK=K<K=K<K;K<K=K>K?K@KAKBKCNKGKFKGKHKIKJKIKJKKKLKMKNKOKPKQKRNKTKUKVKWKXKYNe]�(NKWKVNKTKSKTNKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@NK>K=K<K=K<K;NNK:K;K<K=K>K?K@KAKBKCNKEKFKGKHKIKHKIKJKKKLKMKNKOKPNKRKSKTKUKVKWKXNe]�(NKVKUKTKSKRNKPKOKNKMKLKMNKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K<K;K:K9K:K9K:K;K<K=K>K?K@KAKBKCKDKEKFKGKHKGKHKIKJKKKLKMKNKOKPKQKRNKTKUKVKWNe]�(NKUKTKSKRKQKPKOKNNKLKKNKINKGKFKEKDKCKBKAK@NK>K=K<K;K:K;K:K9K8NK8K9K:K;K<K=K>K?K@KAKBKCKDNNKGKFKGKHKIKJKKKLKMKNKOKPKQKRKSKTKUKVNe]�(NKTKSKRKQKPKOKNKMKLKKKJNKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK9K8K7K8K7K8K9K:K;K<K=K>K?K@KANKCKDKEKFKEKFKGKHKIKJKKKLKMKNKOKPKQKRKSKTKUNe]�(NKSKRKQKPKOKNKMKLKKKJKIKHKGNKEKDKCKBKANK?K>K=K<K;K:K9K8NNK7K6NK6K7K8K9K:K;K<K=K>K?K@KAKBKCNKEKDKEKFKGKHKIKJKKNKOKNKOKPKQKRKSKTNe]�(NKRKQKPKOKNNKNNKJKIKHKGKFKEKDKCKBKAK@K?NK=K<K;NK9K8K7K6K7K6K5K6K5K6K7K8K9K:K;K<K=K>NK@KAKBKCKDKCKDKEKFKGKHKIKJNKNKMKNKOKPKQKRKSNe]�(NKQKPNKNKMKLKMKLKKKJNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K6K5K4K5K4K5K6K7K8K9K:K;K<K=K>K?K@KAKBNKBKCKDKEKFKGKHKIKJNKLKMKNKOKPKQKRNe]�(NKPKOKNKMKLKKKLKMKLKKNKEKDKCKBKCNK?K>K=K<K;NK9NK7NK5K4K5K4K3K4K3K4K5K6K7K8K9K:K;K<K=K>K?K@KAKBKAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQNe]�(NKOKNKMKLKKKJKKKLNNKENKCKBKANK?K>K=K<K;K:NK8K7K6K5NK3K4K3K2K3K2K3K4K5K6K7K8K9K:K;K<K=K>K?K@KAK@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPNe]�(NKNKMKLKKKJKINNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K3K2K1K2K1K2K3K4K5K6K7K8K9K:K;K<K=K>K?K@K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKONe]�(NKMKLKKNKIKHKGKFKENKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K2K1K0K1K0K1K2K3K4K5K6K7K8K9K:K;K<K=K>K?K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNNe]�(NKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0NK0K/NK/K0K1K2K3K4K5K6K7K8K9K:K;K<K=K>K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMNe]�(NKKKJKIKHNKFKENKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4K3NK1K0K/NK/K.K-K.K/K0K1K2K3K4K5K6K7K8K9K:K;K<K=K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLNe]�(NKJNKHKGKFNKDKCKBKCNK?K>K=K<K;K:K9K8NK6K5K4K3K2K1K0K/K.K/K.K-K,K-K.K/K0K1K2K3K4K5K6K7K8K9K:K;K<K;K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKNe]�(NKIKHKGKFKEKDKCKBKANK?K>K=K<K;K:K9K8K7NK5K4K3K2NK0K/NK-K.K-K,K+K,K-K.K/K0K1K2K3K4K5K6K7K8K9K:K;K:K;K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJNe]�(NKHKGKFKEKDKCKBKAK@K?NK=NNK:K9K8K7K6K5K4K3NK1K0K/K.K-K,K-K,K+K*NNNNNNNNNNNNNNNNK9K:K;K<K=K>K?K@NKDKCKDNKFKGKHKINe]�(NKGKFKEKDKCNKAK@K?K>K=K<K;K:K9K8NK6K5K4K3K2NK0K/K.K-K,K+K,K+K*K)NK+K,K-K.K/K0K1K2K3K4K5K6K7K8NK8K9K:K;K<K=K>K?K@NKBKCKDKEKFKGKHNe]�(NKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K1NK/K.K-K,K+K*K+K*K)K(NK*K+K,K-K.K/K0K1K2K3K4K5K6K7NK7K8K9K:K;K<K=K>K?K@KAKBKCKDKEKFKGNe]�(NKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7NK5K4K3K2K1K0K/K.K-K,K+K*K)K*K)K(K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6NK6K7K8K9K:K;K<K=K>K?K@KAKBKCKDKEKFNe]�(NKDKCKBKAK@NNNK<K;K:NK8NK6K5NK3K2K1K0K/K.K-K,K+K*K)K(K)K(K'K&NK*K+K,K-K.K/K0K1K2K3K4K5K6K7NK5K6K7K8K9K:K;K<NK>K?K@KAKBKCKDKENe]�(NKCKBKAK@K?K>NK<K;K:K9K8K7K6K5K4K3K2NK0K/K.K-K,K+K*K)K(K'K(K'K&K%NK+K,K-K.K/K0K1K2K3K4K5K6K7K8NK4K5K6K7K8K9K:K;K<K=K>K?K@KAKBKCKDNe]�(NKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-NK+K*K)K(K'K&K'K&K%K$NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NK3K4K5K6K7K8K9K:K;K<K=K>K?K@NKDKCNe]�(NKANK?K>NK<K;K:NK8K7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K&K%K$K#NNNNNNNNNNNNNNNNK2K3K4K5K6K7K8K9NK;K<K=K>NK@NKBNe]�(NK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K%NK#K"K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1NNK4K5K6K7K8NK:K;K<K=K>K?K@KANe]�(NK?NK=NK;K:K9K8K7NK5K4K3K2K1NK/K.K-K,K+K*K)K(K'NK%NK#NK#K"K!K K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4NK6K7NK9K:K;K<K=K>K?K@Ne]�(NK>K=K<K;K:NK8K7K6NK4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K#K"K!K KK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6NK8K9K:K;K<NK>K?Ne]�(NK=NNK:K9NK7K6K5K4K3NK1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K"K!K KKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2NK4K5K6K7K8K9K:K;K<K=K>Ne]�(NK<K;K:NK8K7K6K5K4K3K2K1K0K/K.K-K,NNK+NK'K&K%K$K#K"K!K K!K NKKKKK K!K"K#K$K%K&K'K(K)K*K+K,NK.K/K0K1K2K3K4NK6K7NNK:K;K<K=Ne]�(NK;K:K9K8K7K6K5K4K3K2K1K0K/K.NK,K+K*K)NNK&K%K$K#K"K!K KK KKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2NK4K5K6K7K8K9K:K;K<Ne]�(NK:K9K8K7K6K5K4K3K2NK0K/K.K-K,K+NK)K(K'K&K%NK#K"K!K KKNKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+NK-K.K/K0K1K2K3K4K5K6K7K8K9K:K;Ne]�(NK9K8K7K6K5NK3K2K1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!K NKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*NK,K-K.K/K0K1K2K3K4NK6K7K8K9K:Ne]�(NK8K7NK5K4K3K2K1K0K/K.K-K,NK*K)NK'K&K%K$K#K"K!K KKKKKKKNKKKKKNKNK!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7K8K9Ne]�(NK7K6K5K4K3K2NK0NK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKNKKK K!K"K#NK%K&NK(K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7K8Ne]�(NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K"NKKKNKKKKKKKKKKKKKNK K!K"K#K$K%K&K'K(NK*K+K,K-NK/K0K1K2K3K4K5K6K7Ne]�(NK5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$NK"K!K NKKKKKNKKKKKNNKNKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6Ne]�(NK4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#NK!K KNKKKKKKKNKKKKKKKNKKKKKK K!K"NK$K%K&K'K(NK*K+NK-K.K/K0K1K2K3K4K5Ne]�(NK3K2K1K0K/K.K-K,NK*K)K(K'NNNNK"K!K KKKKNKKKKKKKKKKKKKNKKKKKKK K!K"K#K$NK(K'K(K)K*K+K,K-K.K/K0K1K2K3K4Ne]�(NK2K1K0K/K.K-NK+NK)K(K'K&K%K$K#K"K!K KNKKKKNKKKNKKKKKKKKKKKKKKNKK K!NK#K$NK&K'K(NK*K+K,K-K.K/K0K1K2K3Ne]�(NK1K0K/K.NK,NK*K)K(K'K&K%K$K#K"K!K NKKKKKKKKKKNKKKKKKKKKKKKNKKKKK K!K"K#K$K%K&K'NK)K*K+K,K-K.K/K0K1K2Ne]�(NK0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKNKKKNKKKKKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1Ne]�(NK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKNKKKKKKKKKKKKKKKKNKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0Ne]�(NK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKNKKKKKKKKKKKKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/Ne]�(NK-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.Ne]�(NK,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKNKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-Ne]�(NK+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKNKKNKKKKKKKKKKKKKNKKNKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,Ne]�(NK*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKNKKKKKKKKKNKKKNKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+Ne]�(NK)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	K
KKKKKKKKKKKNKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*Ne]�(NK(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KNNNNNNNNKKKKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)Ne]�(NK'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKNK	K
KKKKNKKKKKKKKNKKNKKKKK K!K"K#K$K%K&K'K(Ne]�(NK&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKNKK	K
KKKNKKKKKKKKKKKNKKKKKK K!K"K#K$K%K&K'Ne]�(NK%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKKK	K
KKNKKKKKKKKKKKKNKKNKKK K!K"K#K$K%K&Ne]�(NK$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKNKK	K
KKKNKKKKKKKKNKKKKKKKKKKK K!K"K#K$K%Ne]�(NK#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKNK	K
KKKKNKKKKKKKKKKKKKNKKKKKKK K!K"K#K$Ne]�(NK"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKKNK
KKKKKNKKKKKKKKKKNKKKKKKKKKKK K!K"K#Ne]�(NK!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKKKK NNNNNNNK
KKKKKKKKKKKKKKKKKKKKKK K!K"Ne]�(NK"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKKKKKKKKKKK	K
KKKKKKKKKKKKKKKKKKKKKK K!Ne]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�	eliteList�]��Enemies.Goblins��Goblin_Stonewall���a�
messageSys��
MessageSys��Messages���)��}�(�messages�]�(�Player Ready: Kyle��
Game Start�e�retrieveLimit�K�messageLimit�M�ub�healingList�]�h]a�CollisionMap�]�(]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K KKK K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K KK K Ke]�(KK K K K K KK K K K K KKK KK K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K KK K K K KK K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K KK K K K Ke]�(KK K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K KK K K K K K K K K KK K Ke]�(KK K K K K K K K K K KK K K K K K KK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K Ke]�(KK K KK K K K K K K K K KK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K KK K KKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K Ke]�(KK K K K K K K KK K K K K KK K K K K KK KK K K K K K KK K K K K K K K K K K K K KK K K K K K K K K K K K K K K K KK K K K K K Ke]�(KK K KK K K KK K K K K K K K K K K K K K K K K KK K K K K K KKK K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K Ke]�(KK K K K K KK K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K Ke]�(KK K K K K K K K KK K KK KK K K K K K K K KK K K K K K K K K KK K K K K K K K K K K K K KKK K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K KK K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K KK K K K K KK K K K K K K K KKK K KK K K K K K K K K K K K K K KK K K K K K K K K KK K K K K K K K Ke]�(KK K K K K KK KK K K K K K K K K K K K KK K K KK K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K KK K K K K K K K Ke]�(KK K KK K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K KK K K K K K K Ke]�(KK K K K K K K K K K KK K K K K KK K K K K KK KK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K KKK KK K K KK K K K K K KK K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K KKK K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K KK K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K KK K KK K K K K K K K K K K KK K K K K KK K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK KK K K KK K K K KK K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K KK K K K K K K K K KK K K K KK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K KK KKK K K K K K K K KK K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K KK K K KK K K K Ke]�(KK K K K K KK K K K K K K K K K KK K K K K KK K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K KK K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K KK K K K KK K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K Ke]�(KK K K K K KKKK K K KK KK K KK K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K KK K K K K K K K Ke]�(KK K K K K K KK K K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K KK K Ke]�(KK KK K KK K K KK K K K K K K K K K K K K K KK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K KK K K K KK KK Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K KKK K K K K KK K K K K K K K Ke]�(KK KK KK K K K K KK K K K K KK K K K K K K K K KK KK KK K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K Ke]�(KK K K K K KK K K KK K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K KK K Ke]�(KK KKK K KK K K K K KK K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K Ke]�(KK K K KK K K K K K K K K K K K K KKK KK K K K K K K K K K KK K K K K K K K K K K K K K K K K KK K K K K K K KK K KKK K K K Ke]�(KK K K K K K K K K K K K K K KK K K K KKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K Ke]�(KK K K K K K K K K KK K K K K K KK K K K K KK K K K K K KK K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K Ke]�(KK K K K K KK K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K KK K K K K Ke]�(KK K KK K K K K K K K K K KK K KK K K K K K K K K K K K K K K KK K K K K KK KK K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K KK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K KK K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K KK K K K K K KK K K KK K K K K K K K K K K K K KK K K K K K K K K KK K K K KK K K K K K K K K Ke]�(KK K K K K K K K K K K K K K KK K K KK K K KK K K K K KK K K K K KKK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K KK K K KK K K K K K K KK K K K K K K KK K K K K K K K KK K K K K KK K KK K K K K K K K K Ke]�(KK K K K K K K K KK K K K KKKKK K K K K K K KK K K K K K K K K K K K K KK K K K K K K K K K K KK K K K K K K K K K K K K K K Ke]�(KK K K K K K KK KK K K K K K K K K K K KK K K K KK K K KK K K K K K K K K K K K K K KK K K KK K KK K K KK K K K K K K K K K Ke]�(KK K K K KK KK K K K K K K K K K K KK K K K K K K K K K KK K K K K K K K K K K K KK K K K K K K K K K K K KK K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K K K K K K KK K KK K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K KK K K KK K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K KK K KK K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K K K K KK K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K KK K KK K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K KK K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K K K K K K KK K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K K K KK K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKee�	enemyList�]�(j�8  �Goblin_Lancer���j�8  �Goblin_Berserker���j�8  �Goblin_Archer���j�8  �Goblin_Knight���j�8  �Goblin_Grunt���j�8  �Goblin_Thief���e�textWall��Bricks
��	equipList�]�(hh�Iron_Shield���h�Buckler���h�Wooden_Shield���h�	Longsword���h�
Greatsword���h�Bow���h�Spear���h�Dagger���hq�Cloth_Shirt���hshq�Leather_Shirt���hq�Leather_Helm���hq�Iron_Breastplate���hq�	Iron_Helm���hq�Chain_Shirt���hq�
Chain_Helm���eh{h~�djikstra_Player�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NK G�\������G�\�     G�\333333G�[�fffffG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�F������G�F333333G�E������G�E      G�DffffffNe]�(NG�\������G�\�     G�\333333G�[�fffffNNG�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffNG�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      NG�F������G�F333333G�E������G�F333333G�E������NG�DffffffG�C������Ne]�(NG�\�     G�\333333G�[�fffffG�[������G�[L�����NG�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     NNG�X������NG�X      G�W�33333G�WffffffG�W�����G�V�����͕      G�V�     NG�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�E������G�E      G�DffffffG�C������G�C333333Ne]�(NG�\333333G�[�fffffG�[������NG�[      G�Z�33333G�ZffffffG�Z�����NG�Y�     G�Y333333G�X�fffffG�X������G�XL�����NG�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�E      G�DffffffG�C������G�C333333G�B������Ne]�(NG�[�fffffG�[������G�[L�����NG�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      NG�I������G�I333333NG�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������NG�C������G�C333333G�B������G�B      Ne]�(NG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      NG�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffNG�I333333G�H������G�H      NG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�C������G�C333333NG�B      G�AffffffNe]�(NG�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������NG�X      G�W�33333G�WffffffG�W�����G�V������G�V�     NG�U�fffffNG�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������NG�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�C333333G�B������G�B      G�AffffffG�@������Ne]�(NG�[      G�Z�33333NG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333NG�W�����G�V������NG�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffNG�F333333G�E������NG�DffffffG�C������G�C333333G�B������G�B      G�B������G�B      G�AffffffG�@������G�@333333Ne]�(NG�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U������NG�TffffffG�T�����NNG�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      NG�C������G�C333333G�B������G�B      G�AffffffG�B      NG�@������G�@333333G�?333333Ne]�(NG�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�Y�     G�Y333333NG�X      G�W�33333G�WffffffG�W�����G�V������NG�V333333G�U�fffffG�U������G�UL�����G�U      NG�TffffffNG�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����NG�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333NG�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�C333333NG�@������G�AffffffG�@������G�@333333G�?333333G�>      Ne]�(NG�Z�����G�Y������NG�Y333333G�X�fffffG�Y333333NG�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333NG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����NNG�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      NG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      NG�@������G�@333333G�@������G�@333333G�?333333G�>      G�<������Ne]�(NG�Y������G�Y�     G�Y333333G�X�fffffG�X������NG�X      G�W�33333G�WffffffG�W�����G�V������G�W�����NG�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333NG�?333333G�>      G�<������G�;������Ne]�(NG�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffNG�V������G�V�     NG�U�fffffNG�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333NG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333NG�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      NNG�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�?333333G�>      G�<������G�;������G�:ffffffNe]�(NG�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333NG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����NG�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������NG�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�>      G�<������G�;������G�:ffffffG�9333333Ne]�(NG�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����NG�T�33333G�TffffffG�T�����G�S������G�S�     NG�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������NNG�O������G�O333333NG�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333NG�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333NG�>      G�<������G�;������G�<������G�;������G�:ffffffG�9333333G�8      Ne]�(NG�X������G�XL�����G�X      G�W�33333G�WffffffNG�WffffffNG�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffNG�RL�����G�R      G�Q�33333NG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      NG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333NG�<������G�;������G�:ffffffG�;������G�:ffffffG�9333333G�8      G�6������Ne]�(NG�XL�����G�X      NG�WffffffG�W�����G�V������G�W�����G�V������G�V�     G�V333333NG�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffNG�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������NG�:ffffffG�9333333G�:ffffffG�9333333G�8      G�6������G�5������Ne]�(NG�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V������G�W�����G�V������G�V�     NG�T�33333G�TffffffG�T�����G�S������G�T�����NG�R�fffffG�R������G�RL�����G�R      G�Q�33333NG�Q�����NG�P�     NG�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�9333333G�8      G�6������G�5������G�4ffffffNe]�(NG�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�V�     G�V������NNG�T�33333NG�T�����G�S������G�S�     NG�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffNG�P������G�P�     G�P333333G�O������NG�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�8      G�6������G�5������G�4ffffffG�3333333Ne]�(NG�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffNNG�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333NG�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�6������G�5������G�4ffffffG�3333333G�2      Ne]�(NG�W�����G�V������G�V�     NG�U�fffffG�U������G�UL�����G�U      G�T�33333NG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�5������G�4ffffffG�3333333G�2      G�0������Ne]�(NG�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������NG�K������G�K      NG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�4ffffffG�3333333G�2      G�0������G�/333333Ne]�(NG�W�����G�V������G�V�     G�V333333NG�U������G�UL�����NG�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333NG�P�     G�P333333G�O������G�O333333G�N������NG�MffffffG�L������G�L333333NG�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�3333333G�2      G�0������G�/333333G�,������Ne]�(NG�WffffffNG�V������G�V�     G�V333333NG�U������G�UL�����G�U      G�T�33333NG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      NG�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�2      G�0������G�/333333G�,������G�*ffffffNe]�(NG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333NG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333NG�P�     G�P333333G�O������G�O333333NG�N      G�MffffffNG�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�0������G�/333333G�,������G�*ffffffG�(      Ne]�(NG�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����NG�S�     NNG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     NG�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333NNNNNNNNNNNNNNNNG�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333NG�0������G�/333333G�,������NG�,������G�*ffffffG�(      G�%������Ne]�(NG�V�     G�V333333G�U�fffffG�U������G�UL�����NG�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      NG�QffffffG�Q�����G�P������G�P�     G�P333333NG�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������NG�K      G�K������G�L333333G�L������G�MffffffG�N      G�N������G�O333333G�O������G�P333333G�P�     G�P������G�Q�����G�QffffffNG�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������NG�,������G�*ffffffG�(      G�*ffffffG�(      G�%������G�#333333Ne]�(NG�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffNG�P������G�P�     G�P333333G�O������NG�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333NG�JffffffG�K      G�K������G�L333333G�L������G�MffffffG�N      G�N������G�O333333G�O������G�P333333G�P�     G�P������G�Q�����NG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�(      G�%������G�#333333G� ������Ne]�(NG�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����NG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�I333333G�I������G�JffffffG�K      G�K������G�L333333G�L������G�MffffffG�N      G�N������G�O333333G�O������G�P333333G�P�     G�P������NG�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�#333333G�%������G�#333333G� ������G�������Ne]�(NG�V333333G�U�fffffG�U������G�UL�����G�U      NNNG�S������G�S�     G�S333333NG�R������NG�R      G�Q�33333NG�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      NG�JffffffG�K      G�K������G�L333333G�L������G�MffffffG�N      G�N������G�O333333G�O������G�P333333G�P�     G�P������G�Q�����NG�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������NG�(      G�%������G�#333333G� ������G�#333333G� ������G�������G�      Ne]�(NG�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffNG�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������NG�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffNG�K      G�K������G�L333333G�L������G�MffffffG�N      G�N������G�O333333G�O������G�P333333G�P�     G�P������G�Q�����G�QffffffNG�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�#333333G� ������G�������G� ������G�������G�      G�333333Ne]�(NG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������NG�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������NG�K������G�L333333G�L������G�MffffffG�N      G�N������G�O333333G�O������G�P333333G�P�     G�P������G�Q�����G�QffffffG�Q�33333NG�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�#333333G� ������G�������G�      G�������NG�333333G�������Ne]�(NG�UL�����NG�T�33333G�TffffffNG�S������G�S�     G�S333333NG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffNG�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333NNNNNNNNNNNNNNNNG�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffNG� ������G�������G�      G�333333NG�333333NG�333333Ne]�(NG�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������NG�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������NNG�3333333G�2      G�0������G�/333333G�,������NG�������G�      G�333333G�������G�333333G��333333G�       G��333333Ne]�(NG�UL�����NG�T�33333NG�T�����G�S������G�S�     G�S333333G�R�fffffNG�RL�����G�R      G�Q�33333G�QffffffG�Q�����NG�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      NG�I������NG�H������NG�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333NG�0������G�/333333NG� ������G�������G�      G�333333G�������G�333333G��333333G�333333Ne]�(NG�U������G�UL�����G�U      G�T�33333G�TffffffNG�S������G�S�     G�S333333NG�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������NG�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������NG�#333333G� ������G�������G�      G�333333NG�333333G�������Ne]�(NG�U�fffffNNG�TffffffG�T�����NG�S�     G�S333333G�R�fffffG�R������G�RL�����NG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������NG�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333NG�,������G�*ffffffG�(      G�%������G�#333333G� ������G�������G�      G�333333G�������G�333333Ne]�(NG�U������G�UL�����G�U      NG�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333NNG�N������NG�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      NG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffNG�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������NG�(      G�%������NNG�������G�      G�333333G�      Ne]�(NG�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffNG�P������G�P�     G�P333333G�O������NNG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������NG�,������G�*ffffffG�(      G�%������G�#333333G� ������G�������G�      G�������Ne]�(NG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333NG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����NG�O������G�O333333G�N������G�N      G�MffffffNG�L333333G�K������G�K      G�JffffffG�I������G�I333333NG�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333NG�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�#333333G� ������G�������G� ������Ne]�(NG�U�fffffG�U������G�UL�����G�U      G�T�33333NG�T�����G�S������G�S�     G�S333333G�R�fffffNG�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������NG�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffNG�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������NG�(      G�%������G�#333333G� ������G�#333333Ne]�(NG�V333333G�U�fffffNG�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      NG�QffffffG�Q�����NG�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������NG�GffffffG�F������G�F333333G�E������G�E      NG�C������NG�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�#333333G�%������Ne]�(NG�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffNG�S������NG�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������NG�DffffffG�C������G�C333333G�B������G�B      G�AffffffNG�@333333G�?333333NG�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�%������G�(      Ne]�(NG�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333NG�Q�����G�P������G�P�     G�P333333G�O������G�O333333NG�N      G�MffffffG�L������NG�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffNG�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������NG�:ffffffG�9333333G�8      G�6������NG�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�(      G�*ffffffNe]�(NG�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������NG�R      G�Q�33333G�QffffffNG�P������G�P�     G�P333333NG�O333333G�N������G�N      G�MffffffG�N      NG�K������G�K      G�JffffffG�I������G�I333333NNG�GffffffNG�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�*ffffffG�,������Ne]�(NG�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333NG�Q�����G�P������G�P�     NG�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333NG�K      G�JffffffG�I������G�I333333G�H������G�H      G�H������NG�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      NG�@������G�@333333G�?333333G�>      G�<������NG�:ffffffG�9333333NG�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�,������G�/333333Ne]�(NG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      NG�TffffffG�T�����G�S������G�S�     NNNNG�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333NG�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�I333333NG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������NG�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�/333333G�0������Ne]�(NG�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffNG�UL�����NG�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333NG�Q�����G�P������G�P�     G�P������NG�O333333G�N������G�N      NG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      NG�C������G�C333333G�B������NG�AffffffG�B      NG�?333333G�>      G�<������NG�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�0������G�2      Ne]�(NG�W�33333G�WffffffG�W�����G�V������NG�V333333NG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������NG�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������NG�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������NG�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      NG�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�2      G�3333333Ne]�(NG�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333NG�O333333G�N������G�N      NG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�3333333G�4ffffffNe]�(NG�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     NG�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������NG�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�4ffffffG�5������Ne]�(NG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����NG�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�5������G�6������Ne]�(NG�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�6������G�8      Ne]�(NG�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333NG�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�8      G�9333333Ne]�(NG�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      NG�QffffffG�Q�����NG�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������NG�H������G�H      NG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�9333333G�:ffffffNe]�(NG�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     NG�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      NG�I������G�I333333G�H������NG�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�:ffffffG�;������Ne]�(NG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������NG�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�;������G�<������Ne]�(NG�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������NNNNNNNNG�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�<������G�>      Ne]�(NG�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����NG�R�fffffG�S333333G�S�     G�S������G�T�����G�TffffffNG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������NG�GffffffG�F������NG�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�>      G�?333333Ne]�(NG�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffNG�R������G�R�fffffG�S333333G�S�     G�S������G�T�����NG�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffNG�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�?333333G�@333333Ne]�(NG�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�R      G�RL�����G�R������G�R�fffffG�S333333G�S�     G�S������NG�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�H������NG�F333333G�E������NG�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�@333333G�@������Ne]�(NG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      NG�R������G�R�fffffG�S333333G�S�     G�S������G�T�����NG�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffNG�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�@������G�AffffffNe]�(NG�[�fffffG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����NG�R�fffffG�S333333G�S�     G�S������G�T�����G�TffffffNG�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      NG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�AffffffG�B      Ne]�(NG�\333333G�[�fffffG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������NG�S333333G�S�     G�S������G�T�����G�TffffffG�T�33333NG�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffNG�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�B      G�B������Ne]�(NG�\�     G�\333333G�[�fffffG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�S333333NNNNNNNG�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�B������G�C333333Ne]�(NG�\������G�\�     G�\333333G�[�fffffG�[������G�[L�����G�[      G�Z�33333G�ZffffffG�Z�����G�Y������G�Y�     G�Y333333G�X�fffffG�X������G�XL�����G�X      G�W�33333G�WffffffG�W�����G�V������G�V�     G�V333333G�U�fffffG�U������G�UL�����G�U      G�T�33333G�TffffffG�T�����G�S������G�S�     G�S333333G�R�fffffG�R������G�RL�����G�R      G�Q�33333G�QffffffG�Q�����G�P������G�P�     G�P333333G�O������G�O333333G�N������G�N      G�MffffffG�L������G�L333333G�K������G�K      G�JffffffG�I������G�I333333G�H������G�H      G�GffffffG�F������G�F333333G�E������G�E      G�DffffffG�C������G�C333333G�C������Ne]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�levelManager��LevelManager�j�9  ��)��}�(�	gameState�h)��}�(hK#h�hKKhKh	h�	levelList�j�9  �MessageHandler�j�8  �height�K�gameVersion��0.1.0��console��tdl��Console���)��KYKE]�(K K K K ��K K K ����KKK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KLK�K�K���K K K ����KEK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KRK�K�K���K K K ����KPK�K�K���K K K ����KAK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KWK�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KGK�K�K���K K K ����KPK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KxK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KaK�K�K���K K K ����KoK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����KFK�K�K���K K K ����K K K K ��K K K ����KvK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KnK�K�K���K K K ����KwK�K�K���K K K ����KmK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KmK�K�K���K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KwK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K0K�K�K���K K K ����K K K K ��K K K ����KhK�K�K���K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K:K�K�K���K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KSK�K�K���K K K ����KrK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KPK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KtK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K1K�K�K���K K K ����K2K�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����KRK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K9K�K�K���K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KrK�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KBK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KtK�K�K���K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KFK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����e(K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KKK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K��      K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����e(K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����e(K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K@KKYK���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����e(K K�K�K���K K K ����K K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K �����       K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����e(K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����e��b�xConst�K,ubj�9  ]�h�aj�8  j�8  �nextSeed�M�M�cursor�K ub�inSeed�M��	textSpace��ground, covered in leaves
��maze�]�(]�(�T�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  �.�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �~�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  h"j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �x�j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  haj��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �#�jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �D�j��  j��  j��  j��  j��  j��  j��  j��  �=�j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  h"j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �X�j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �S�j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  haj��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jс  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j΁  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  haj��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j́  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jс  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  h"j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  haj��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  jс  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  �E�jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  ee�djikstra_Player_Away�jQ9  �SeesMap�]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK KK K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K Ke]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK KKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK KKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K KKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKK K K K K KKKK e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K KKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K ee�args�]�(KKe�SeenMap�]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK KK K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K Ke]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK KKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K �       K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK KKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K KKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKK K K K K KKKK e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K KKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K eej�9  j�9  �djikstra_Stairs_Up�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NKaK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K&K%K$K#K"Ne]�(NK`K_K^K]NNKZKYKXKWKVKUKTKSKRKQKPKOKNNKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K%K$NK"K!Ne]�(NK_K^K]K\K[NKYKXKWKVKUNNKRNKPKOKNKMKLKKNKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K$K#K"K!K Ne]�(NK^K]K\NKZKYKXKWNKUKTKSKRKQNKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K#K"K!K KNe]�(NK]K\K[NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-NK+K*NK(K'K&K%K$K#K"K!NK!K KKNe]�(NK\K[KZKYKXKWKVKUKTKSKRKQKPNKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,NK*K)K(NK&K%K$K#K"K!K K!K NKKNe]�(NK[KZKYKXKWKVKUKTKSKRNKPKOKNKMKLKKNKINKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K!K KK KKKKNe]�(NKZKYNKWKVKUKTKSKRKQKPKONKMKLNKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$NK"K!K KKKKKKKNe]�(NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKHNKDKCNNK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#NK!K KKKKNKKKNe]�(NKXKWKVKUKTKUKTNKPKOKNKMKLNKJKIKHKGKFNKDNKBKAK@K?K>K=NK;K:K9K8K7K6K5K4K3K2K1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!K KK NKKKKKKNe]�(NKWKVNKTKSKTNKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@NK>K=K<K;K:K9NNK6K5K4K3K2K1K0K/K.K-NK+K*K)K(K'K&K%K$K#K"K!K KKNKKKKKKKNe]�(NKVKUKTKSKRNKPKOKNKMKLKMNKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKNKKKKNe]�(NKUKTKSKRKQKPKOKNNKLKKNKINKGKFKEKDKCKBKAK@NK>K=K<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+K*K)K(NNK%K$K#K"K!K KKKKKKKKKKKKNe]�(NKTKSKRKQKPKOKNKMKLKKKJNKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4K3K2K1K0K/K.K-K,K+K*K)NK'K&K%K$K#K"K!K KKKKKKKKKKKKKNe]�(NKSKRKQKPKOKNKMKLKKKJKIKHKGNKEKDKCKBKANK?K>K=K<K;K:K9K8NNK5K4NK2K1K0K/K.K-K,K+K*K)K(K'K&K%NK#K"K!K KKKKKNKKKKKKKKNe]�(NKRKQKPKOKNNKNNKJKIKHKGKFKEKDKCKBKAK@K?NK=K<K;NK9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K KKKKKKNKKKKKKKKNe]�(NKQKPNKNKMKLKMKLKKKJNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"NK KKKKKKKKNKKKKKKKNe]�(NKPKOKNKMKLKKKLKMKLKKNKEKDKCKBKCNK?K>K=K<K;NK9NK7NK5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKNe]�(NKOKNKMKLKKKJKKKLNNKENKCKBKANK?K>K=K<K;K:NK8K7K6K5NK3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKNe]�(NKNKMKLKKKJKINNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKNe]�(NKMKLKKNKIKHKGKFKENKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKNe]�(NKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0NK.K-NK+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKNe]�(NKMKLKKKJNKHKGNKEKDKCKBKAK@K?K>K=K<K;NK7K6K5K4K3NK1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKNe]�(NKNNKLKKKJNKHKGKFKENKCKBKAK@K?K>K=K<NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKNe]�(NKMKLKKKJKIKHKGKFKENKCKBKAK@K?K>K=K<K;NK7K6K5K4NK2K1NK-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKK
Ne]�(NKLKKKJKIKHKGKFKEKDKCNKANNK>K=K<K;K:K9K8K7NK3K2K1K0K/K.K-K,K+K*NNNNNNNNNNNNNNNNKKKKKKKKNKKKNKKK
K	Ne]�(NKKKJKIKHKGNKEKDKCKBKAK@K?K>K=K<NK:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+NK-K.K/K0K1K2K3K4K5K6K7K8K9K:NKKKKKKKKKNKKK
KK
K	KNe]�(NKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK8K7K6K5NK3K2K1K0K/K.K-K,K+K*NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NKKKKKKKKKKKK
K	K
K	KKNe]�(NKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=NK9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7K8NKKKKKKKKKKK
K	KK	KKKNe]�(NKJKIKHKGKFNNNKBKAK@NK>NK<K;NK7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NKKKKKKKKNK
K	KKKKKKNe]�(NKIKHKGKFKEKDNKBKAK@K?K>K=K<K;K:K9K8NK4K3K2K1K0K/K.K-K,K+K*K)K(K'NK-K.K/K0K1K2K3K4K5K6K7K8K9K:NKKKKKKKKK
K	KKKKKKKNe]�(NKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3NK/K.K-K,K+K*K)K(K'K&NK.K/K0K1K2K3K4K5K6K7K8K9K:K;NKKKKKKKK
K	KKKKKNKKNe]�(NKGNKEKDNKBKAK@NK>K=K<K;K:K9K8K7K6K5K4K3K2K1NK-K,K+K*K)K(K'K&K%NNNNNNNNNNNNNNNNKKKKKKKKNKKKKNKNKNe]�(NKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)NK%K$K#K"K!K KKKKKKKKKKKKKNNKKKKKNKKKKKKK KNe]�(NKGNKENKCKBKAK@K?NK=K<K;K:K9NK5K4K3K2K1K0K/K.K-NK+NK)NK'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKNKKNKKKKKKKKNe]�(NKHKGKFKEKDNKBKAK@NK<K;K:K9K8K7K6K5K4K3NK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKNKKKKKNKKNe]�(NKINNKDKCNKAK@K?K>K=NK9K8K7K6K5K4K3K2K1K0NK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKNKKK
K	KKKKKKKNe]�(NKHKGKFNKBKAK@K?K>K=K<K;K:K9K8K7K6NNK3NK1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K KKKKKKKKKKNKKKKKKKNK
K	NNKKKKNe]�(NKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK8K7K6K5NNK0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKNKKK
K	KKKKKNe]�(NKHKGKFKEKDKCKBKAK@NK>K=K<K;K:K9NK5K4K3K2K1NK/K.K-K,K+K*NK(K'K&K%K$K#K"K!K KKKKKKKKKKKNKKKKKKKKKK
K	KKKKNe]�(NKIKHKGKFKENKCKBKAK@K?NK;K:K9K8K7K6K5K4K3K2K1K0K/K.NK,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKNKKKKKKKKKNK
K	KKKNe]�(NKJKINKEKDKCKBKAK@K?K>K=K<NK:K9NK7K6K5K4K3K2K1K0K/K.K-K,K+K*K)NK'K&K%K$K#NK!NKKKKKKKKKKKKKKKKKKKKKK
K	KK	Ne]�(NKIKHKGKFKEKDNKBNK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$NK"K!K KKKNKKNKKKKKKKKKKKKKKK
K	K
Ne]�(NKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;NK9K8K7K6K5K4NK2K1K0NK.K-K,K+K*K)K(K'K&K%K$K#K"NK KKKKKKKKNKKKKNKKKKKKKK
KNe]�(NKKKJKIKHKGKFKEKDKCKBKAK@K?K>NK<K;K:NK8K7K6NK4K3K2K1K2NK.K-K,K+K*NNK'NK%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKNe]�(NKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;NK9K8K7NK5K4K3K2K1K0K/NK-K,K+K*K)K(K)NK%K$K#K"K!K KKNKKKKKNKKNKKKKKKKKKNe]�(NKMKLKKKJKIKHKGKFNKDKCKBKANNNNK<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+K*K)K*NK&K%K$K#K"K!K KKKKNKKKKKKKKKKKKKKKNe]�(NKNKMKLKKKJKINKGNKEKDKCKBKAK@K?K>K=K<K;NK9K8K7K8NK4K3K2NK0K/K.K-K,K+K*K)K(K'K&K%K$K#NK!K KNKKNKKKNKKKKKKKKKKNe]�(NKOKNKMKLNKJNKHKGKFKEKDKCKBKAK@K?K>NK<K;K:K9K8K7K6K5K4K3NK1K0K/K.K-K,K+K*K)K(K'K&NK$K#K"K!K KKKKKKKNKKKKKKKKKKNe]�(NKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2NK0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKNe]�(NKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7NK5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&NK$K#K"K!K KKKKKKKKKKKKKKKKNe]�(NKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKNe]�(NKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKNe]�(NKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*NK(K'K&K%K$K#K"K!K KKKKKKKKKKKKKNe]�(NKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NK:K9NK7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(NK&K%K$K#K"K!K KKKKKKKKKKKKNe]�(NKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7NK5K4K3K2K1K0K/K.K-NK+K*K)NK'K&K%K$K#K"K!K KKKKKKKKKKKNe]�(NKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K!K KKKKKKKKKKNe]�(NKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8NNNNNNNNK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKNe]�(NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK?K@KAKBKCKDNK0K/K.K-K,K+K*K)NK'K&NK$K#K"K!K KKKKKKKKNe]�(NKZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK>K?K@KAKBKCNK1K0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K KKKKKKKNe]�(NK[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K<K=K>K?K@KAKBNK2K1K0K/K.K-K,K+K*K)K(K)NK%K$NK"K!K KKKKKKNe]�(NK\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NK>K?K@KAKBKCNK3K2K1K0K/K.K-K,NK*K)K(K'K&K%K$K#K"K!K KKKKKNe]�(NK]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=NK?K@KAKBKCKDNK4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K KKKKNe]�(NK^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>NK@KAKBKCKDKENK5K4K3K2K1K0K/K.K-K,NK*K)K(K'K&K%K$K#K"K!K KKKNe]�(NK_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K@NNNNNNNK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KK Ne]�(NK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K K!Ne]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�stairsUp�]�(K"KAe�itemList�]�(h]h[�Bundle_Of_Arrows���h[�	Time_Bomb���h[�Scroll_of_Fireball���h[�Scroll_of_Lightning_Bolt���hj39  j59  j79  j99  j;9  j=9  j?9  jA9  jC9  hsjE9  jG9  jI9  jK9  jM9  jO9  ej  }�(K h})��}�(h�Kh�K h!h"h�h�j  K'h&�Item�h|j=9  )��}�(h{jڂ  hKhKhKhhhhh�h�hKh �h!h"h#Kh$�h%Kh&�Bow�h(�ububKh})��}�(h�Kh�Kh!j��  h�h�j  K#h&�Enemy�h|j'9  )��}�(hK
hK hj=9  )��}�(hKhKhKhhhhh�h�hKh �h!h"h#Kh$�h%Kh&j߂  h(�ubhKh)�h*��isAfraid��h+Kh,�h!j��  h7K	hKh8K hK hphs)��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&hvhhwub�	cowardice�G?�      hfKhNN�lastPlayerMap�Nhn]�hPKdhRKh&�Goblin Archer�hTK hY]�hMK hg]�h]�(K�KKe�lastPlayerLoc�NhjK �
dropChance�K(�
stealthVal�K �necklace�NhO�hmNhxKhy��hearingDist�Kh{j��  �armor�jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&�Leather Shirt�h�armor�ub�
alliesList�]�(j��  h})��}�(h�Kh�Kh!j��  h�h�j  K'h&j�  h|j)9  )��}�(hKhK hj99  )��}�(hKhKhKhhh�1H�h�h�hKh �h!h"h#Kh$�h%Kh&�	Longsword�h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjK9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&�	Iron Helm�hhwubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&�Goblin Knight�hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j��  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j��  hj��  ubj��  ]�(j��  j��  e�leftHand�j79  )��}�(hKhKhhhj�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&�Wooden Shield�hK ub�blocking��h%Kububej�  Nj�  �h%KububKj��  Kh})��}�(h�Kh�Kh!j��  h�h�j  K8h&j�  h|j+9  )��}�(hK	hK hj99  )��}�(hKhKhKhhhj�  h�h�hKh �h!h"h#Kh$�h%Kh&j�  h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hhh&�Leather Helm�hhwubj�  G?��Q�hfKhNNj�  Nhn]�hPKdhRKh&�Goblin Grunt�hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j��  hj��  ubj��  ]�(j�  h})��}�(h�Kh�Kh!j��  h�h�j  K6h&j�  h|j%9  )��}�(hKhK hj;9  )��}�(hKhKhKhhhhh�h�hKh �h!h"h#Kh$�h%Kh&�
Greatsword�h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hhh&j�  hhwubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&�Goblin Berserker�hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j$�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j��  hj��  ubj��  ]�(j�  j$�  ej�  Nj�  �h%Kububej�  Nj�  �h%KububKh})��}�(h�Kh�Kh!hah�h�j  K5h&�Health�h|h])��}�(h`Kh�h(�h!hah{j4�  hhh&hbhhcububKj$�  Kh})��}�(h�Kh�Kh!j��  h�h�j  K(h&j�  h|j'9  )��}�(hK
hK hj=9  )��}�(hKhKhKhhhhh�h�hKh �h!h"h#Kh$�h%Kh&j߂  h(�ubhKh)�h*�j�  �h+Kh,�h!j��  h7KhKh8K hK hphs)��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&hvhhwubj�  G?�      hfKhNNj�  Nhn]�hPKdhRKh&j�  hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j9�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j��  hj��  ubj��  ]�(j9�  h})��}�(h�Kh�Kh!j��  h�h�j  K+h&j�  h|j#9  )��}�(hK	hK hj?9  )��}�(hKhKhKhhhhh�h�hKh �h!h"h#Kh$�h%Kh&�Spear�h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hhh&j�  hhwubj�  G?�������hfKhNNj�  Nhn]�hPKdhRKh&�Goblin Lancer�hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{jG�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j��  hj��  ubj��  ]�(j9�  jG�  h})��}�(h�Kh�K
h!j��  h�h�j  K#h&j�  h|j%9  )��}�(hKhK hj;9  )��}�(hKhKhKhhhhh�h�hKh �h!h"h#Kh$�h%Kh&j*�  h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hhh&j�  hhwubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&j.�  hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{jW�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j��  hj��  ubj��  ]�(j9�  jW�  ej�  Nj�  �h%Kububh})��}�(h�Kh�Kh!jс  h�h�j  K.h&j�  h|j�8  )��}�(hKhK hh�Mace���)��}�(hKhKhKhhhj�  h�h�hKh �h!h"h#Kh$�h%Kh&�Mace�h(�ubhKh)�h*�j�  �h+K h,�h!jс  h7K	hKh8K hK hpjK9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j�  hhwubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&�Goblin Stonewall�hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{je�  j��  jI9  )��}�(h�h(�hKh!h"h#K7h8K2h$�hhh&�Iron Breastplate�hj��  ubj��  ]�(jG�  je�  ej�  j39  )��}�(hKhKhhhj�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&�Iron Shield�hK ubj�  �h%Kububej�  j59  )��}�(hKhKhhh�0H�h�h�h(�h �h!h"h#Kh8Kh$�h%K h&�Buckler�hK ubj�  �h%KububjW�  je�  ej�  Nj�  �h%KububKjG�  Kh})��}�(h�Kh�Kh!j΁  h�h�j  K+h&�Chest�h|�Features.Features��Chest���)��}�(h{j�  hY]�(jM9  )��}�(h�h(�hKh!h"h#K#h8K#h$�hhh&�Chain Shirt�hj��  ubjA9  )��}�(hKhKhKhhhj�  h�h�hKh �h!h"h#Kh$�h%Kh&�Dagger�h(�ubj79  )��}�(hKhKhhhj�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&j�  hK ubh[�
Gold_Coins���)��}�(h��coins�Kh(�h!�$�h]�(K�K�Keh&�
Gold Coins�hhcubeh!j΁  h]�(KQKOKeh&j��  ububK	h})��}�(h�Kh�K	h!h"h�h�j  K(h&j܂  h|j79  )��}�(h{j��  hKhKhhhj�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&j�  hK ububK
jW�  Kje�  Kh})��}�(h�K"h�Kh!jՁ  h�h�j  KAh&�	Stairs Up�h|�Features.Stairs��StairUp���)��}�(h{j��  h�K"h�J����h�h�j  KA�moveCost�Kh&�Stairs�h|NububKh~Kh})��}�(h�K5h�Kh!hah�h�j  K=h&j6�  h|h])��}�(h`Kh�h(�h!hah{j��  hhh&hbhhcububKh})��}�(h�K7h�Kh!jс  h�h�j  K=h&j�  h|j�8  )��}�(hKhK hjj�  )��}�(hKhKhKhhhj�  h�h�hKh �h!h"h#Kh$�h%Kh&jm�  h(�ubhKh)�h*�j�  �h+K h,�h!jс  h7KhKh8K hK hpjK9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j�  hhwubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&jq�  hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j��  j��  jI9  )��}�(h�h(�hKh!h"h#K7h8K2h$�hhh&jv�  hj��  ubj��  ]�j�  j39  )��}�(hKhKhhhj�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&jz�  hK ubj�  �h%KububKh})��}�(h�K7h�Kh!j��  h�h�j  K@h&j�  h|j%9  )��}�(hKhK hj;9  )��}�(hKhKhKhhhhh�h�hKh �h!h"h#Kh$�h%Kh&j*�  h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hhh&j�  hhwubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&j.�  hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j��  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j��  hj��  ubj��  ]�j�  Nj�  �h%KububKh})��}�(h�K;h�Kh!j΁  h�h�j  Kh&j��  h|j��  )��}�(h{jɃ  hY]�(j39  )��}�(hKhKhhhj�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&jz�  hK ubj39  )��}�(hKhKhhhj�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&jz�  hK ubhs)��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&hvhhwubj��  )��}�(h�j��  Kh(�h!j��  hj��  h&j��  hhcubeh!j΁  hj��  h&j��  ububKh})��}�(h�K<h�Kh!j��  h�h�j  Kh&j�  h|j%9  )��}�(hKhK hj;9  )��}�(hKhKhKhhhhh�h�hKh �h!h"h#Kh$�h%Kh&j*�  h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hhh&j�  hhwubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&j.�  hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{jփ  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j��  hj��  ubj��  ]�j�  Nj�  �h%KububKh})��}�(h�K=h�Kh!j��  h�h�j  Kh&j�  h|j+9  )��}�(hK	hK hj99  )��}�(hKhKhKhhhj�  h�h�hKh �h!h"h#Kh$�h%Kh&j�  h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hhh&j�  hhwubj�  G?��Q�hfKhNNj�  Nhn]�hPKdhRKh&j�  hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j��  hj��  ubj��  ]�j�  Nj�  �h%KububKh})��}�(h�K=h�Kh!j��  h�h�j  Kh&j�  h|j'9  )��}�(hK
hK hj=9  )��}�(hKhKhKhhhhh�h�hKh �h!h"h#Kh$�h%Kh&j߂  h(�ubhKh)�h*�j�  �h+Kh,�h!j��  h7KhKh8K hK hphs)��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&hvhhwubj�  G?�      hfKhNNj�  Nhn]�hPKdhRKh&j�  hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j��  hj��  ubj��  ]�j�  Nj�  �h%KububKh})��}�(h�K=h�Kh!hah�h�j  Kh&j6�  h|h])��}�(h`Kh�h(�h!hah{j �  hhh&hbhhcububKh})��}�(h�K>h�Kh!j��  h�h�j  Kh&j�  h|j'9  )��}�(hK
hK hj=9  )��}�(hKhKhKhhhhh�h�hKh �h!h"h#Kh$�h%Kh&j߂  h(�ubhKh)�h*�j�  �h+Kh,�h!j��  h7KhKh8K hK hphs)��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&hvhhwubj�  G?�      hfKhNNj�  Nhn]�hPKdhRKh&j�  hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j��  hj��  ubj��  ]�j�  Nj�  �h%KububKh})��}�(h�K>h�Kh!jс  h�h�j  Kh&j�  h|j�8  )��}�(hKhK hjj�  )��}�(hKhKhKhhhj�  h�h�hKh �h!h"h#Kh$�h%Kh&jm�  h(�ubhKh)�h*�j�  �h+K h,�h!jс  h7KhKh8K hK hpjK9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j�  hhwubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&jq�  hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j�  j��  jI9  )��}�(h�h(�hKh!h"h#K7h8K2h$�hhh&jv�  hj��  ubj��  ]�j�  j39  )��}�(hKhKhhhj�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&jz�  hK ubj�  �h%KububKh})��}�(h�K?h�Kh!h"h�h�j  Kh&j܂  h|j59  )��}�(h{j"�  hKhKhhhj}�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&j~�  hK ububKh})��}�(h�K?h�Kh!hah�h�j  K'h&j6�  h|h])��}�(h`Kh�h(�h!hah{j&�  hhh&hbhhcububKh})��}�(h�K@h�Kh!jс  h�h�j  K$h&j�  h|j�8  )��}�(hKhK hjj�  )��}�(hKhKhKhhhj�  h�h�hKh �h!h"h#Kh$�h%Kh&jm�  h(�ubhKh)�h*�j�  �h+K h,�h!jс  h7K	hKh8K hK hpjK9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j�  hhwubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&jq�  hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j*�  j��  jI9  )��}�(h�h(�hKh!h"h#K7h8K2h$�hhh&jv�  hj��  ubj��  ]�j�  j39  )��}�(hKhKhhhj�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&jz�  hK ubj�  �h%KububKh})��}�(h�K@h�Kh!j��  h�h�j  K%h&j�  h|j%9  )��}�(hKhK hj;9  )��}�(hKhKhKhhhhh�h�hKh �h!h"h#Kh$�h%Kh&j*�  h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hhh&j�  hhwubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&j.�  hTK hY]�hMK hg]�hj��  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j:�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&j��  hj��  ubj��  ]�j�  Nj�  �h%KububKh})��}�(h�KAh�Kh!j��  h�h�j  K"h&�Stairs Down�h|j��  �	StairDown���)��}�(h{jH�  h|Nh�J����h�h�h�KAj��  Kh&j��  j  K"ububu�consumeList�]�(h]j҂  jԂ  jւ  j؂  eh&�
1B: Forest��djikstra_Player_Adj�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K%K$K#K"K!Ne]�(NK_K^K]K\NNKYKXKWKVKUKTKSKRKQKPKOKNKMNKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$K#K$K#NK!K Ne]�(NK^K]K\K[KZNKXKWKVKUKTNNKQNKOKNKMKLKKKJNKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K#K"K!K KNe]�(NK]K\K[NKYKXKWKVNKTKSKRKQKPNKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K"K!K KKNe]�(NK\K[KZNKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,NK*K)NK'K&K%K$K#K"K!K NK KKKNe]�(NK[KZKYKXKWKVKUKTKSKRKQKPKONKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(K'NK%K$K#K"K!K KK KNKKNe]�(NKZKYKXKWKVKUKTKSKRKQNKOKNKMKLKKKJNKHNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*NK(K'K&K%K$K#K"K!K KKKKKKKNe]�(NKYKXNKVKUKTKSKRKQKPKOKNNKLKKNKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&NK$K#NK!K KKKKKKKKNe]�(NKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKGNKCKBNNK?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"NK KKKKKNKKKNe]�(NKWKVKUKTKSKTKSNKOKNKMKLKKNKIKHKGKFKENKCNKAK@K?K>K=K<NK:K9K8K7K6K5K4K3K2K1K0K/K.NK,K+K*K)K(K'K&K%K$K#K"K!K KKKNKKKKKKNe]�(NKVKUNKSKRKSNKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?NK=K<K;K:K9K8NNK5K4K3K2K1K0K/K.K-K,NK*K)K(K'K&K%K$K#K"K!K KKKNKKKKKKKNe]�(NKUKTKSKRKQNKOKNKMKLKKKLNKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKNKKKKNe]�(NKTKSKRKQKPKOKNKMNKKKJNKHNKFKEKDKCKBKAK@K?NK=K<K;K:K9K8K7K6K5NK3K2K1K0K/K.K-K,K+K*K)K(K'NNK$K#K"K!K KKKKKKKKKKKKKNe]�(NKSKRKQKPKOKNKMKLKKKJKINKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K KKKKKKKKKKKKKKNe]�(NKRKQKPKOKNKMKLKKKJKIKHKGKFNKDKCKBKAK@NK>K=K<K;K:K9K8K7NNK4K3NK1K0K/K.K-K,K+K*K)K(K'K&K%K$NK"K!K KKKKKKNKKKKKKKKNe]�(NKQKPKOKNKMNKMNKIKHKGKFKEKDKCKBKAK@K?K>NK<K;K:NK8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K KKKKKKKNKKKKKKKKNe]�(NKPKONKMKLKKKLKKKJKINKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!NKKKKKKKKKNKKKKKKKNe]�(NKOKNKMKLKKKJKKKLKKKJNKDKCKBKAKBNK>K=K<K;K:NK8NK6NK4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKNe]�(NKNKMKLKKKJKIKJKKNNKDNKBKAK@NK>K=K<K;K:K9NK7K6K5K4NK2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKNe]�(NKMKLKKKJKIKHNNKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5NK3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKNe]�(NKLKKKJNKHKGKFKEKDNKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKNe]�(NKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/NK-K,NK*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKNe]�(NKLKKKJKINKGKFNKDKCKBKAK@K?K>K=K<K;K:NK6K5K4K3K2NK0K/K.NK,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKNe]�(NKMNKKKJKINKGKFKEKDNKBKAK@K?K>K=K<K;NK5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKK
Ne]�(NKLKKKJKIKHKGKFKEKDNKBKAK@K?K>K=K<K;K:NK6K5K4K3NK1K0NK,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKK
K	Ne]�(NKKKJKIKHKGKFKEKDKCKBNK@NNK=K<K;K:K9K8K7K6NK2K1K0K/K.K-K,K+K*K)NNNNNNNNNNNNNNNNKKKKKKKKNKKKNKK
K	KNe]�(NKJKIKHKGKFNKDKCKBKAK@K?K>K=K<K;NK9K8K7K6K5NK3K2K1K0K/K.K-K,K+K*NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NKKKKKKKKKNKK
K	K
K	KKNe]�(NKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4NK2K1K0K/K.K-K,K+K*K)NK+K,K-K.K/K0K1K2K3K4K5K6K7K8NKKKKKKKKKKK
K	KK	KKKNe]�(NKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NK8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7NKKKKKKKKKK
K	KKKKKKNe]�(NKIKHKGKFKENNNKAK@K?NK=NK;K:NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK+K,K-K.K/K0K1K2K3K4K5K6K7K8NKKKKKKKKNK	KKKKKKKNe]�(NKHKGKFKEKDKCNKAK@K?K>K=K<K;K:K9K8K7NK3K2K1K0K/K.K-K,K+K*K)K(K'K&NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NKKKKKKKK
K	KKKKKKKKNe]�(NKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2NK.K-K,K+K*K)K(K'K&K%NK-K.K/K0K1K2K3K4K5K6K7K8K9K:NKKKKKKK
K	KKKKKKNKKNe]�(NKFNKDKCNKAK@K?NK=K<K;K:K9K8K7K6K5K4K3K2K1K0NK,K+K*K)K(K'K&K%K$NNNNNNNNNNNNNNNNKKKKKKKK
NKKKKNKK KNe]�(NKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK$K#K"K!K KKKKKKKKKKKKKKNNKKKKKNKKKKKK KK Ne]�(NKFNKDNKBKAK@K?K>NK<K;K:K9K8NK4K3K2K1K0K/K.K-K,NK*NK(NK&K%K$K#K"K!K KKKKKKKKKKKKKKKKKNKKNKKKKKKK KNe]�(NKGKFKEKDKCNKAK@K?NK;K:K9K8K7K6K5K4K3K2NK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKNKKKKKNKKNe]�(NKHNNKCKBNK@K?K>K=K<NK8K7K6K5K4K3K2K1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKNKK
K	KKKKKKKKNe]�(NKGKFKENKAK@K?K>K=K<K;K:K9K8K7K6K5NNK2NK0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K KKKKKKKKKKKNKKKKKKKNK	KNNKKKKNe]�(NKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4NNK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKNKK
K	KKKKKKNe]�(NKGKFKEKDKCKBKAK@K?NK=K<K;K:K9K8NK4K3K2K1K0NK.K-K,K+K*K)NK'K&K%K$K#K"K!K KKKKKKKKKKKKNKKKKKKKKK
K	KKKKKNe]�(NKHKGKFKEKDNKBKAK@K?K>NK:K9K8K7K6K5K4K3K2K1K0K/K.K-NK+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKNKKKKKKKKKNK	KKKKNe]�(NKIKHNKDKCKBKAK@K?K>K=K<K;NK9K8NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"NK NKKKKKKKKKKKKKKKKKKKKK
K	KKKNe]�(NKHKGKFKEKDKCNKANK?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#NK!K KKKKNKKNKKKKKKKKKKKKKK
K	KK	Ne]�(NKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK8K7K6K5K4K3NK1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!NKKKKKKKKKNKKKKNKKKKKKK
K	K
Ne]�(NKJKIKHKGKFKEKDKCKBKAK@K?K>K=NK;K:K9NK7K6K5NK3K2K1K0K1NK-K,K+K*K)NNK&NK$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
KNe]�(NKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK8K7K6NK4K3K2K1K0K/K.NK,K+K*K)K(K'K(NK$K#K"K!K KKKNKKKKKNKKNKKKKKKKKKNe]�(NKLKKKJKIKHKGKFKENKCKBKAK@NNNNK;K:K9K8K7K6K5NK3K2K1K0K/K.K-K,K+K*K)K(K)NK%K$K#K"K!K KKKKKNKKKKKKKKKKKKKKKNe]�(NKMKLKKKJKIKHNKFNKDKCKBKAK@K?K>K=K<K;K:NK8K7K6K7NK3K2K1NK/K.K-K,K+K*K)K(K'K&K%K$K#K"NK KKNKKNKKKNKKKKKKKKKKNe]�(NKNKMKLKKNKINKGKFKEKDKCKBKAK@K?K>K=NK;K:K9K8K7K6K5K4K3K2NK0K/K.K-K,K+K*K)K(K'K&K%NK#K"K!K KKKKKKKKNKKKKKKKKKKNe]�(NKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5NK3K2K1NK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKNe]�(NKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%NK#K"K!K KKKKKKKKKKKKKKKKKNe]�(NKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKNe]�(NKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKNe]�(NKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)NK'K&K%K$K#K"K!K KKKKKKKKKKKKKKNe]�(NKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;NK9K8NK6K5K4K3K2K1K0K/K.K-K,K+K*NK(K'NK%K$K#K"K!K KKKKKKKKKKKKKNe]�(NKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,NK*K)K(NK&K%K$K#K"K!K KKKKKKKKKKKKNe]�(NKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*NK(K'K&K%K$K#K"K!K KKKKKKKKKKKNe]�(NKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7NNNNNNNNK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKNe]�(NKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8NK>K?K@KAKBKCNK/K.K-K,K+K*K)K(NK&K%NK#K"K!K KKKKKKKKKNe]�(NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK=K>K?K@KAKBNK0K/K.K-K,K+K*K)K(K'K&NK$K#K"K!K KKKKKKKKNe]�(NKZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K;K<K=K>K?K@KANK1K0K/K.K-K,K+K*K)K(K'K(NK$K#NK!K KKKKKKKNe]�(NK[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;NK=K>K?K@KAKBNK2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K!K KKKKKKNe]�(NK\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NK>K?K@KAKBKCNK3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K KKKKKNe]�(NK]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=NK?K@KAKBKCKDNK4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K!K KKKKNe]�(NK^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K?NNNNNNNK5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKNe]�(NK_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KK Ne]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�cLevel�Kubj  KAh&�Player�h|hubj��  jC9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hhh&�Cloth Shirt�hj��  ubj�  h�Tome���)��}�(hK hKhKhhhj}�  h�h�hKh �h!h"h#Kh$�h%K h&�Tome�h(�ubj�  �j�  Nubj�9  j�9  )��}�(j�9  hj�9  ]�h�)��}�(h�]�(h�h�h�eh	h)��}�(hKhK hh)��}�(hKhKhKh]�(K�K�K�eh�2H�h�h�hKh �h!h"h#Kh$�h%Kh&�Staff�h(�ubhKh)�h*�h+K h,�h!h-h.}�(h0K h1K h2K h3K h4K h5K h6K uh7K hKh8K hK h9Nh:Kh%Kh;K�h<}�(h0h@h1hBh2hDh3hFh4hHh5hJh6hLuhMK hNNhO�hPKdhQG?�      hRK�h&�Kyle�hTK hUhXhY]�(h])��}�(h`Kh�h(�h!hahj��  h&�
Green Herb�h�
consumable�ubh])��}�(h`Kh�h(�h!hahj��  h&j��  hj��  ubehfKhg]�h]�(KKYK�ehjK hkNhlK hmNhn]�hphs)��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&�	Cloth Hat�h�helmet�ubhxK�hy�hzK h{h})��}�(h�K$h�Kh!h-h�j��  j  K?h&�Player�h|j��  ubj��  jC9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&�Cloth Shirt�h�armor�ubj�  j��  )��}�(hK hKhKhj��  h�0H�h�h�hKh �h!h"h#Kh$�h%K h&�Tome�h(�ubj�  �j�  Nubh�]�(]�(K#K>e]�(K"K=e]�(K!K<e]�(K K;e]�(KK:e]�(KK9e]�(KK8e]�(KK7e]�(K#K@e]�(K"KAe]�(K!KBe]�(K KCe]�(K#K>e]�(K"K=e]�(K!K<e]�(K K;e]�(KK:e]�(KK9e]�(KK8e]�(KK7e]�(K#K@e]�(K"KAe]�(K!KBe]�(K KCe]�(K#K>e]�(K"K=e]�(K!K<e]�(K!K;e]�(K K:e]�(KK9e]�(KK8e]�(KK7e]�(K#K@e]�(K"KAe]�(K"KBe]�(K!KCe]�(K#K>e]�(K"K=e]�(K"K<e]�(K!K;e]�(K K:e]�(KK9e]�(KK8e]�(KK7e]�(K#K@e]�(K#KAe]�(K"KBe]�(K!KCe]�(K#K>e]�(K#K=e]�(K"K<e]�(K!K;e]�(K!K:e]�(K#K@e]�(K#KAe]�(K"KBe]�(K!KCe]�(K#K>e]�(K#K=e]�(K"K<e]�(K"K;e]�(K!K:e]�(K#K@e]�(K#KAe]�(K"KBe]�(K"KCe]�(K#K>e]�(K#K=e]�(K"K<e]�(K"K;e]�(K!K:e]�(K$K@e]�(K$K>e]�(K#K=e]�(K#K<e]�(K"K;e]�(K"K:e]�(K$K@e]�(K$K>e]�(K#K=e]�(K#K<e]�(K#K;e]�(K"K:e]�(K$K@e]�(K$K>e]�(K#K=e]�(K#K<e]�(K#K;e]�(K#K:e]�(K$K@e]�(K$K>e]�(K$K=e]�(K#K<e]�(K#K;e]�(K#K:e]�(K$K@e]�(K$K>e]�(K$K=e]�(K$K<e]�(K$K;e]�(K$K:e]�(K$K@e]�(K$K>e]�(K$K=e]�(K$K<e]�(K$K;e]�(K$K:e]�(K$K@e]�(K$K>e]�(K$K=e]�(K$K<e]�(K$K;e]�(K$K:e]�(K$K@e]�(K$K>e]�(K$K=e]�(K%K<e]�(K%K;e]�(K%K:e]�(K%K9e]�(K%K8e]�(K%K7e]�(K$K@e]�(K$K>e]�(K%K=e]�(K%K<e]�(K%K;e]�(K%K:e]�(K&K9e]�(K&K8e]�(K&K7e]�(K$K@e]�(K$K>e]�(K%K=e]�(K%K<e]�(K%K;e]�(K&K:e]�(K$K@e]�(K$K>e]�(K%K=e]�(K%K<e]�(K&K;e]�(K&K:e]�(K$K@e]�(K%K>e]�(K%K=e]�(K&K<e]�(K&K;e]�(K'K:e]�(K'K9e]�(K$K@e]�(K%K>e]�(K%K=e]�(K&K<e]�(K&K;e]�(K'K:e]�(K(K9e]�(K(K8e]�(K)K7e]�(K%K@e]�(K%KAe]�(K&KBe]�(K&KCe]�(K%K>e]�(K%K=e]�(K&K<e]�(K'K;e]�(K'K:e]�(K(K9e]�(K)K8e]�(K)K7e]�(K%K@e]�(K%KAe]�(K&KBe]�(K'KCe]�(K%K>e]�(K&K=e]�(K%K@e]�(K%KAe]�(K&KBe]�(K'KCe]�(K%K>e]�(K&K=e]�(K%K@e]�(K&KAe]�(K&KBe]�(K'KCe]�(K%K>e]�(K&K=e]�(K%K@e]�(K&KAe]�(K'KBe]�(K(KCe]�(K%K>e]�(K&K=e]�(K%K@e]�(K&KAe]�(K'KBe]�(K(KCe]�(K#K>e]�(K"K=e]�(K!K<e]�(K K;e]�(KK:e]�(KK9e]�(KK8e]�(KK7e]�(K%K>e]�(K&K=e]�(K#K>e]�(K"K=e]�(K!K<e]�(K K;e]�(KK:e]�(KK9e]�(KK9e]�(KK8e]�(K%K>e]�(K&K=e]�(K#K>e]�(K"K=e]�(K!K<e]�(K K<e]�(KK;e]�(KK:e]�(K%K>e]�(K&K=e]�(K#K>e]�(K"K=e]�(K!K=e]�(K K<e]�(KK;e]�(KK:e]�(K%K>e]�(K&K>e]�(K#K>e]�(K"K>e]�(K!K=e]�(K K<e]�(KK<e]�(KK;e]�(KK:e]�(KK:e]�(K%K>e]�(K&K>e]�(K#K>e]�(K"K>e]�(K!K=e]�(K K=e]�(KK<e]�(KK;e]�(KK;e]�(KK:e]�(K%K>e]�(K&K>e]�(K#K>e]�(K"K>e]�(K!K=e]�(K K=e]�(KK<e]�(KK<e]�(KK;e]�(KK;e]�(K%K?e]�(K&K>e]�(K#K?e]�(K"K>e]�(K!K>e]�(K K=e]�(KK=e]�(KK<e]�(KK<e]�(KK<e]�(K%K?e]�(K&K>e]�(K#K?e]�(K"K>e]�(K!K>e]�(K K>e]�(KK=e]�(KK=e]�(KK=e]�(KK<e]�(K%K?e]�(K&K>e]�(K#K?e]�(K"K>e]�(K!K>e]�(K K>e]�(KK>e]�(KK=e]�(KK=e]�(KK=e]�(K%K?e]�(K&K?e]�(K'K>e]�(K(K>e]�(K)K>e]�(K*K>e]�(K+K=e]�(K,K=e]�(K#K?e]�(K"K?e]�(K!K>e]�(K K>e]�(KK>e]�(KK>e]�(KK>e]�(KK>e]�(K%K?e]�(K&K?e]�(K'K?e]�(K(K>e]�(K)K>e]�(K*K>e]�(K+K>e]�(K,K>e]�(K#K?e]�(K"K?e]�(K!K?e]�(K%K?e]�(K&K?e]�(K'K?e]�(K(K?e]�(K)K?e]�(K*K?e]�(K+K>e]�(K,K>e]�(K#K?e]�(K"K?e]�(K!K?e]�(K%K?e]�(K&K?e]�(K'K?e]�(K(K?e]�(K)K?e]�(K*K?e]�(K+K?e]�(K,K?e]�(K#K?e]�(K"K?e]�(K!K?e]�(K%K?e]�(K&K?e]�(K'K?e]�(K(K?e]�(K)K?e]�(K*K?e]�(K+K@e]�(K,K@e]�(K#K?e]�(K"K?e]�(K!K@e]�(K K@e]�(K%K?e]�(K&K?e]�(K'K?e]�(K(K@e]�(K)K@e]�(K*K@e]�(K+K@e]�(K,K@e]�(K#K?e]�(K"K@e]�(K!K@e]�(K K@e]�(K%K?e]�(K&K?e]�(K'K@e]�(K(K@e]�(K)K@e]�(K*K@e]�(K+KAe]�(K,KAe]�(K#K?e]�(K"K@e]�(K!K@e]�(K K@e]�(K%K?e]�(K&K@e]�(K'K@e]�(K(K@e]�(K)KAe]�(K*KAe]�(K+KAe]�(K,KBe]�(K#K?e]�(K"K@e]�(K!K@e]�(K KAe]�(KKAe]�(KKBe]�(KKBe]�(KKBe]�(K%K?e]�(K&K@e]�(K'K@e]�(K(KAe]�(K)KAe]�(K*KAe]�(K+KBe]�(K,KBe]�(K#K@e]�(K"K@e]�(K!KAe]�(K%K?e]�(K&K@e]�(K'K@e]�(K(KAe]�(K)KAe]�(K*KBe]�(K+KBe]�(K,KCe]�(K#K@e]�(K"K@e]�(K!KAe]�(K%K@e]�(K&K@e]�(K'KAe]�(K(KAe]�(K)KBe]�(K*KBe]�(K+KCe]�(K#K@e]�(K"K@e]�(K!KAe]�(K%K@e]�(K&K@e]�(K'KAe]�(K(KBe]�(K)KBe]�(K*KCe]�(K#K@e]�(K"KAe]�(K!KAe]�(K%K@e]�(K&K@e]�(K'KAe]�(K(KBe]�(K)KCe]�(K#K@e]�(K"KAe]�(K!KBe]�(K KBe]�(KKCe]�(K%K@e]�(K&KAe]�(K'KAe]�(K(KBe]�(K)KCe]�(K#K@e]�(K"KAe]�(K!KBe]�(K KCe]�(K%K@e]�(K&KAe]�(K'KBe]�(K(KCe]�(K#K@e]�(K"KAe]�(K!KBe]�(K KCe]�(K%K@e]�(K&KAe]�(K'KBe]�(K(KCeej  ]�(KAK"ej  }�(K }�(K j	  )��}�(h�K j  ]�h�j��  j  K ubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubK	j	  )��}�(h�K j  ]�h�j��  j  K	ubK
j	  )��}�(h�K j  ]�h�j��  j  K
ubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubK j	  )��}�(h�K j  ]�h�j��  j  K ubK!j	  )��}�(h�K j  ]�h�j��  j  K!ubK"j	  )��}�(h�K j  ]�h�j��  j  K"ubK#j	  )��}�(h�K j  ]�h�j��  j  K#ubK$j	  )��}�(h�K j  ]�h�j��  j  K$ubK%j	  )��}�(h�K j  ]�h�j��  j  K%ubK&j	  )��}�(h�K j  ]�h�j��  j  K&ubK'j	  )��}�(h�K j  ]�h�j��  j  K'ubK(j	  )��}�(h�K j  ]�h�j��  j  K(ubK)j	  )��}�(h�K j  ]�h�j��  j  K)ubK*j	  )��}�(h�K j  ]�h�j��  j  K*ubK+j	  )��}�(h�K j  ]�h�j��  j  K+ubK,j	  )��}�(h�K j  ]�h�j��  j  K,ubK-j	  )��}�(h�K j  ]�h�j��  j  K-ubK.j	  )��}�(h�K j  ]�h�j��  j  K.ubK/j	  )��}�(h�K j  ]�h�j��  j  K/ubK0j	  )��}�(h�K j  ]�h�j��  j  K0ubK1j	  )��}�(h�K j  ]�h�j��  j  K1ubK2j	  )��}�(h�K j  ]�h�j��  j  K2ubK3j	  )��}�(h�K j  ]�h�j��  j  K3ubK4j	  )��}�(h�K j  ]�h�j��  j  K4ubK5j	  )��}�(h�K j  ]�h�j��  j  K5ubK6j	  )��}�(h�K j  ]�h�j��  j  K6ubK7j	  )��}�(h�K j  ]�h�j��  j  K7ubK8j	  )��}�(h�K j  ]�h�j��  j  K8ubK9j	  )��}�(h�K j  ]�h�j��  j  K9ubK:j	  )��}�(h�K j  ]�h�j��  j  K:ubK;j	  )��}�(h�K j  ]�h�j��  j  K;ubK<j	  )��}�(h�K j  ]�h�j��  j  K<ubK=j	  )��}�(h�K j  ]�h�j��  j  K=ubK>j	  )��}�(h�K j  ]�h�j��  j  K>ubK?j	  )��}�(h�K j  ]�h�j��  j  K?ubK@j	  )��}�(h�K j  ]�h�j��  j  K@ubKAj	  )��}�(h�K j  ]�h�j��  j  KAubKBj	  )��}�(h�K j  ]�h�j��  j  KBubKCj	  )��}�(h�K j  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�K ah�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�Kah�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�Kah�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK	}�(K j	  )��}�(h�K	j  ]�h�j��  j  K ubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubK	j	  )��}�(h�K	j  ]�h�j��  j  K	ubK
j	  )��}�(h�K	j  ]�h�j��  j  K
ubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubKj	  )��}�(h�K	j  ]�h�j��  j  KubK j	  )��}�(h�K	j  ]�h�j��  j  K ubK!j	  )��}�(h�K	j  ]�h�j��  j  K!ubK"j	  )��}�(h�K	j  ]�h�j��  j  K"ubK#j	  )��}�(h�K	j  ]�h�j��  j  K#ubK$j	  )��}�(h�K	j  ]�h�j��  j  K$ubK%j	  )��}�(h�K	j  ]�h�j��  j  K%ubK&j	  )��}�(h�K	j  ]�h�j��  j  K&ubK'j	  )��}�(h�K	j  ]�h�j��  j  K'ubK(j	  )��}�(h�K	j  ]�h�j��  j  K(ubK)j	  )��}�(h�K	j  ]�h�j��  j  K)ubK*j	  )��}�(h�K	j  ]�h�j��  j  K*ubK+j	  )��}�(h�K	j  ]�h�j��  j  K+ubK,j	  )��}�(h�K	j  ]�h�j��  j  K,ubK-j	  )��}�(h�K	j  ]�h�j��  j  K-ubK.j	  )��}�(h�K	j  ]�h�j��  j  K.ubK/j	  )��}�(h�K	j  ]�h�j��  j  K/ubK0j	  )��}�(h�K	j  ]�h�j��  j  K0ubK1j	  )��}�(h�K	j  ]�h�j��  j  K1ubK2j	  )��}�(h�K	j  ]�h�j��  j  K2ubK3j	  )��}�(h�K	j  ]�h�j��  j  K3ubK4j	  )��}�(h�K	j  ]�h�j��  j  K4ubK5j	  )��}�(h�K	j  ]�h�j��  j  K5ubK6j	  )��}�(h�K	j  ]�h�j��  j  K6ubK7j	  )��}�(h�K	j  ]�h�j��  j  K7ubK8j	  )��}�(h�K	j  ]�h�j��  j  K8ubK9j	  )��}�(h�K	j  ]�h�j��  j  K9ubK:j	  )��}�(h�K	j  ]�h�j��  j  K:ubK;j	  )��}�(h�K	j  ]�h�j��  j  K;ubK<j	  )��}�(h�K	j  ]�h�j��  j  K<ubK=j	  )��}�(h�K	j  ]�h�j��  j  K=ubK>j	  )��}�(h�K	j  ]�h�j��  j  K>ubK?j	  )��}�(h�K	j  ]�h�j��  j  K?ubK@j	  )��}�(h�K	j  ]�h�j��  j  K@ubKAj	  )��}�(h�K	j  ]�h�j��  j  KAubKBj	  )��}�(h�K	j  ]�h�j��  j  KBubKCj	  )��}�(h�K	j  ]�h�j��  j  KCubuK
}�(K j	  )��}�(h�K
j  ]�h�j��  j  K ubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubK	j	  )���       }�(h�K
j  ]�h�j��  j  K	ubK
j	  )��}�(h�K
j  ]�h�j��  j  K
ubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubKj	  )��}�(h�K
j  ]�h�j��  j  KubK j	  )��}�(h�K
j  ]�h�j��  j  K ubK!j	  )��}�(h�K
j  ]�h�j��  j  K!ubK"j	  )��}�(h�K
j  ]�h�j��  j  K"ubK#j	  )��}�(h�K
j  ]�h�j��  j  K#ubK$j	  )��}�(h�K
j  ]�h�j��  j  K$ubK%j	  )��}�(h�K
j  ]�h�j��  j  K%ubK&j	  )��}�(h�K
j  ]�h�j��  j  K&ubK'j	  )��}�(h�K
j  ]�h�j��  j  K'ubK(j	  )��}�(h�K
j  ]�h�j��  j  K(ubK)j	  )��}�(h�K
j  ]�h�j��  j  K)ubK*j	  )��}�(h�K
j  ]�h�j��  j  K*ubK+j	  )��}�(h�K
j  ]�h�j��  j  K+ubK,j	  )��}�(h�K
j  ]�h�j��  j  K,ubK-j	  )��}�(h�K
j  ]�h�j��  j  K-ubK.j	  )��}�(h�K
j  ]�h�j��  j  K.ubK/j	  )��}�(h�K
j  ]�h�j��  j  K/ubK0j	  )��}�(h�K
j  ]�h�j��  j  K0ubK1j	  )��}�(h�K
j  ]�h�j��  j  K1ubK2j	  )��}�(h�K
j  ]�h�j��  j  K2ubK3j	  )��}�(h�K
j  ]�h�j��  j  K3ubK4j	  )��}�(h�K
j  ]�h�j��  j  K4ubK5j	  )��}�(h�K
j  ]�h�j��  j  K5ubK6j	  )��}�(h�K
j  ]�h�j��  j  K6ubK7j	  )��}�(h�K
j  ]�h�j��  j  K7ubK8j	  )��}�(h�K
j  ]�h�j��  j  K8ubK9j	  )��}�(h�K
j  ]�h�j��  j  K9ubK:j	  )��}�(h�K
j  ]�h�j��  j  K:ubK;j	  )��}�(h�K
j  ]�h�j��  j  K;ubK<j	  )��}�(h�K
j  ]�h�j��  j  K<ubK=j	  )��}�(h�K
j  ]�h�j��  j  K=ubK>j	  )��}�(h�K
j  ]�h�j��  j  K>ubK?j	  )��}�(h�K
j  ]�h�j��  j  K?ubK@j	  )��}�(h�K
j  ]�h�j��  j  K@ubKAj	  )��}�(h�K
j  ]�h�j��  j  KAubKBj	  )��}�(h�K
j  ]�h�j��  j  KBubKCj	  )��}�(h�K
j  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�Kah�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�Kah�j��  j  K5ubK6j	  )��}�(h�Kj  ]�Kah�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�Kah�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�Kah�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�Kah�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�h�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�K	ah�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�h�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK}�(K j	  )��}�(h�Kj  ]�h�j��  j  K ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK	j	  )��}�(h�Kj  ]�h�j��  j  K	ubK
j	  )��}�(h�Kj  ]�h�j��  j  K
ubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubKj	  )��}�(h�Kj  ]�h�j��  j  KubK j	  )��}�(h�Kj  ]�h�j��  j  K ubK!j	  )��}�(h�Kj  ]�h�j��  j  K!ubK"j	  )��}�(h�Kj  ]�h�j��  j  K"ubK#j	  )��}�(h�Kj  ]�K
ah�j��  j  K#ubK$j	  )��}�(h�Kj  ]�h�j��  j  K$ubK%j	  )��}�(h�Kj  ]�h�j��  j  K%ubK&j	  )��}�(h�Kj  ]�h�j��  j  K&ubK'j	  )��}�(h�Kj  ]�h�j��  j  K'ubK(j	  )��}�(h�Kj  ]�h�j��  j  K(ubK)j	  )��}�(h�Kj  ]�h�j��  j  K)ubK*j	  )��}�(h�Kj  ]�h�j��  j  K*ubK+j	  )��}�(h�Kj  ]�h�j��  j  K+ubK,j	  )��}�(h�Kj  ]�h�j��  j  K,ubK-j	  )��}�(h�Kj  ]�h�j��  j  K-ubK.j	  )��}�(h�Kj  ]�Kah�j��  j  K.ubK/j	  )��}�(h�Kj  ]�h�j��  j  K/ubK0j	  )��}�(h�Kj  ]�h�j��  j  K0ubK1j	  )��}�(h�Kj  ]�h�j��  j  K1ubK2j	  )��}�(h�Kj  ]�h�j��  j  K2ubK3j	  )��}�(h�Kj  ]�h�j��  j  K3ubK4j	  )��}�(h�Kj  ]�h�j��  j  K4ubK5j	  )��}�(h�Kj  ]�h�j��  j  K5ubK6j	  )��}�(h�Kj  ]�h�j��  j  K6ubK7j	  )��}�(h�Kj  ]�h�j��  j  K7ubK8j	  )��}�(h�Kj  ]�h�j��  j  K8ubK9j	  )��}�(h�Kj  ]�h�j��  j  K9ubK:j	  )��}�(h�Kj  ]�h�j��  j  K:ubK;j	  )��}�(h�Kj  ]�h�j��  j  K;ubK<j	  )��}�(h�Kj  ]�h�j��  j  K<ubK=j	  )��}�(h�Kj  ]�h�j��  j  K=ubK>j	  )��}�(h�Kj  ]�h�j��  j  K>ubK?j	  )��}�(h�Kj  ]�h�j��  j  K?ubK@j	  )��}�(h�Kj  ]�h�j��  j  K@ubKAj	  )��}�(h�Kj  ]�h�j��  j  KAubKBj	  )��}�(h�Kj  ]�h�j��  j  KBubKCj	  )��}�(h�Kj  ]�h�j��  j  KCubuK }�(K j	  )��}�(h�K j  ]�h�j��  j  K ubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubK	j	  )��}�(h�K j  ]�h�j��  j  K	ubK
j	  )��}�(h�K j  ]�h�j��  j  K
ubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubKj	  )��}�(h�K j  ]�h�j��  j  KubK j	  )��}�(h�K j  ]�h�j��  j  K ubK!j	  )��}�(h�K j  ]�h�j��  j  K!ubK"j	  )��}�(h�K j  ]�h�j��  j  K"ubK#j	  )��}�(h�K j  ]�h�j��  j  K#ubK$j	  )��}�(h�K j  ]�h�j��  j  K$ubK%j	  )��}�(h�K j  ]�h�j��  j  K%ubK&j	  )��}�(h�K j  ]�h�j��  j  K&ubK'j	  )��}�(h�K j  ]�h�j��  j  K'ubK(j	  )��}�(h�K j  ]�h�j��  j  K(ubK)j	  )��}�(h�K j  ]�h�j��  j  K)ubK*j	  )��}�(h�K j  ]�h�j��  j  K*ubK+j	  )��}�(h�K j  ]�h�j��  j  K+ubK,j	  )��}�(h�K j  ]�h�j��  j  K,ubK-j	  )��}�(h�K j  ]�h�j��  j  K-ubK.j	  )��}�(h�K j  ]�h�j��  j  K.ubK/j	  )��}�(h�K j  ]�h�j��  j  K/ubK0j	  )��}�(h�K j  ]�h�j��  j  K0ubK1j	  )��}�(h�K j  ]�h�j��  j  K1ubK2j	  )��}�(h�K j  ]�h�j��  j  K2ubK3j	  )��}�(h�K j  ]�h�j��  j  K3ubK4j	  )��}�(h�K j  ]�h�j��  j  K4ubK5j	  )��}�(h�K j  ]�h�j��  j  K5ubK6j	  )��}�(h�K j  ]�h�j��  j  K6ubK7j	  )��}�(h�K j  ]�h�j��  j  K7ubK8j	  )��}�(h�K j  ]�h�j��  j  K8ubK9j	  )��}�(h�K j  ]�h�j��  j  K9ubK:j	  )��}�(h�K j  ]�h�j��  j  K:ubK;j	  )��}�(h�K j  ]�h�j��  j  K;ubK<j	  )��}�(h�K j  ]�h�j��  j  K<ubK=j	  )��}�(h�K j  ]�h�j��  j  K=ubK>j	  )��}�(h�K j  ]�h�j��  j  K>ubK?j	  )��}�(h�K j  ]�h�j��  j  K?ubK@j	  )��}�(h�K j  ]�h�j��  j  K@ubKAj	  )��}�(h�K j  ]�h�j��  j  KAubKBj	  )��}�(h�K j  ]�h�j��  j  KBubKCj	  )��}�(h�K j  ]�h�j��  j  KCubuK!}�(K j	  )��}�(h�K!j  ]�h�j��  j  K ubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubK	j	  )��}�(h�K!j  ]�h�j��  j  K	ubK
j	  )��}�(h�K!j  ]�h�j��  j  K
ubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubKj	  )��}�(h�K!j  ]�h�j��  j  KubK j	  )��}�(h�K!j  ]�h�j��  j  K ubK!j	  )��}�(h�K!j  ]�h�j��  j  K!ubK"j	  )��}�(h�K!j  ]�h�j��  j  K"ubK#j	  )��}�(h�K!j  ]�h�j��  j  K#ubK$j	  )��}�(h�K!j  ]�h�j��  j  K$ubK%j	  )��}�(h�K!j  ]�h�j��  j  K%ubK&j	  )��}�(h�K!j  ]�h�j��  j  K&ubK'j	  )��}�(h�K!j  ]�h�j��  j  K'ubK(j	  )��}�(h�K!j  ]�h�j��  j  K(ubK)j	  )��}�(h�K!j  ]�h�j��  j  K)ubK*j	  )��}�(h�K!j  ]�h�j��  j  K*ubK+j	  )��}�(h�K!j  ]�h�j��  j  K+ubK,j	  )��}�(h�K!j  ]�h�j��  j  K,ubK-j	  )��}�(h�K!j  ]�h�j��  j  K-ubK.j	  )��}�(h�K!j  ]�h�j��  j  K.ubK/j	  )��}�(h�K!j  ]�h�j��  j  K/ubK0j	  )��}�(h�K!j  ]�h�j��  j  K0ubK1j	  )��}�(h�K!j  ]�h�j��  j  K1ubK2j	  )��}�(h�K!j  ]�h�j��  j  K2ubK3j	  )��}�(h�K!j  ]�h�j��  j  K3ubK4j	  )��}�(h�K!j  ]�h�j��  j  K4ubK5j	  )��}�(h�K!j  ]�h�j��  j  K5ubK6j	  )��}�(h�K!j  ]�h�j��  j  K6ubK7j	  )��}�(h�K!j  ]�h�j��  j  K7ubK8j	  )��}�(h�K!j  ]�h�j��  j  K8ubK9j	  )��}�(h�K!j  ]�h�j��  j  K9ubK:j	  )��}�(h�K!j  ]�h�j��  j  K:ubK;j	  )��}�(h�K!j  ]�h�j��  j  K;ubK<j	  )��}�(h�K!j  ]�h�j��  j  K<ubK=j	  )��}�(h�K!j  ]�h�j��  j  K=ubK>j	  )��}�(h�K!j  ]�h�j��  j  K>ubK?j	  )��}�(h�K!j  ]�h�j��  j  K?ubK@j	  )��}�(h�K!j  ]�h�j��  j  K@ubKAj	  )��}�(h�K!j  ]�h�j��  j  KAubKBj	  )��}�(h�K!j  ]�h�j��  j  KBubKCj	  )��}�(h�K!j  ]�h�j��  j  KCubuK"}�(K j	  )��}�(h�K"j  ]�h�j��  j  K ubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubK	j	  )��}�(h�K"j  ]�h�j��  j  K	ubK
j	  )��}�(h�K"j  ]�h�j��  j  K
ubKj	  )��}�(h��      K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubKj	  )��}�(h�K"j  ]�h�j��  j  KubK j	  )��}�(h�K"j  ]�h�j��  j  K ubK!j	  )��}�(h�K"j  ]�h�j��  j  K!ubK"j	  )��}�(h�K"j  ]�h�j��  j  K"ubK#j	  )��}�(h�K"j  ]�h�j��  j  K#ubK$j	  )��}�(h�K"j  ]�h�j��  j  K$ubK%j	  )��}�(h�K"j  ]�h�j��  j  K%ubK&j	  )��}�(h�K"j  ]�h�j��  j  K&ubK'j	  )��}�(h�K"j  ]�h�j��  j  K'ubK(j	  )��}�(h�K"j  ]�h�j��  j  K(ubK)j	  )��}�(h�K"j  ]�h�j��  j  K)ubK*j	  )��}�(h�K"j  ]�h�j��  j  K*ubK+j	  )��}�(h�K"j  ]�h�j��  j  K+ubK,j	  )��}�(h�K"j  ]�h�j��  j  K,ubK-j	  )��}�(h�K"j  ]�h�j��  j  K-ubK.j	  )��}�(h�K"j  ]�h�j��  j  K.ubK/j	  )��}�(h�K"j  ]�h�j��  j  K/ubK0j	  )��}�(h�K"j  ]�h�j��  j  K0ubK1j	  )��}�(h�K"j  ]�h�j��  j  K1ubK2j	  )��}�(h�K"j  ]�h�j��  j  K2ubK3j	  )��}�(h�K"j  ]�h�j��  j  K3ubK4j	  )��}�(h�K"j  ]�h�j��  j  K4ubK5j	  )��}�(h�K"j  ]�h�j��  j  K5ubK6j	  )��}�(h�K"j  ]�h�j��  j  K6ubK7j	  )��}�(h�K"j  ]�h�j��  j  K7ubK8j	  )��}�(h�K"j  ]�h�j��  j  K8ubK9j	  )��}�(h�K"j  ]�h�j��  j  K9ubK:j	  )��}�(h�K"j  ]�h�j��  j  K:ubK;j	  )��}�(h�K"j  ]�h�j��  j  K;ubK<j	  )��}�(h�K"j  ]�h�j��  j  K<ubK=j	  )��}�(h�K"j  ]�h�j��  j  K=ubK>j	  )��}�(h�K"j  ]�h�j��  j  K>ubK?j	  )��}�(h�K"j  ]�h�j��  j  K?ubK@j	  )��}�(h�K"j  ]�h�j��  j  K@ubKAj	  )��}�(h�K"j  ]�Kah�j��  j  KAubKBj	  )��}�(h�K"j  ]�h�j��  j  KBubKCj	  )��}�(h�K"j  ]�h�j��  j  KCubuK#}�(K j	  )��}�(h�K#j  ]�h�j��  j  K ubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubK	j	  )��}�(h�K#j  ]�h�j��  j  K	ubK
j	  )��}�(h�K#j  ]�h�j��  j  K
ubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubKj	  )��}�(h�K#j  ]�h�j��  j  KubK j	  )��}�(h�K#j  ]�h�j��  j  K ubK!j	  )��}�(h�K#j  ]�h�j��  j  K!ubK"j	  )��}�(h�K#j  ]�h�j��  j  K"ubK#j	  )��}�(h�K#j  ]�h�j��  j  K#ubK$j	  )��}�(h�K#j  ]�h�j��  j  K$ubK%j	  )��}�(h�K#j  ]�h�j��  j  K%ubK&j	  )��}�(h�K#j  ]�h�j��  j  K&ubK'j	  )��}�(h�K#j  ]�h�j��  j  K'ubK(j	  )��}�(h�K#j  ]�h�j��  j  K(ubK)j	  )��}�(h�K#j  ]�h�j��  j  K)ubK*j	  )��}�(h�K#j  ]�h�j��  j  K*ubK+j	  )��}�(h�K#j  ]�h�j��  j  K+ubK,j	  )��}�(h�K#j  ]�h�j��  j  K,ubK-j	  )��}�(h�K#j  ]�h�j��  j  K-ubK.j	  )��}�(h�K#j  ]�h�j��  j  K.ubK/j	  )��}�(h�K#j  ]�h�j��  j  K/ubK0j	  )��}�(h�K#j  ]�h�j��  j  K0ubK1j	  )��}�(h�K#j  ]�h�j��  j  K1ubK2j	  )��}�(h�K#j  ]�h�j��  j  K2ubK3j	  )��}�(h�K#j  ]�h�j��  j  K3ubK4j	  )��}�(h�K#j  ]�h�j��  j  K4ubK5j	  )��}�(h�K#j  ]�h�j��  j  K5ubK6j	  )��}�(h�K#j  ]�h�j��  j  K6ubK7j	  )��}�(h�K#j  ]�h�j��  j  K7ubK8j	  )��}�(h�K#j  ]�h�j��  j  K8ubK9j	  )��}�(h�K#j  ]�h�j��  j  K9ubK:j	  )��}�(h�K#j  ]�h�j��  j  K:ubK;j	  )��}�(h�K#j  ]�h�j��  j  K;ubK<j	  )��}�(h�K#j  ]�h�j��  j  K<ubK=j	  )��}�(h�K#j  ]�h�j��  j  K=ubK>j	  )��}�(h�K#j  ]�h�j��  j  K>ubK?j	  )��}�(h�K#j  ]�h�j��  j  K?ubK@j	  )��}�(h�K#j  ]�h�j��  j  K@ubKAj	  )��}�(h�K#j  ]�h�j��  j  KAubKBj	  )��}�(h�K#j  ]�h�j��  j  KBubKCj	  )��}�(h�K#j  ]�h�j��  j  KCubuK$}�(K j	  )��}�(h�K$j  ]�h�j��  j  K ubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubK	j	  )��}�(h�K$j  ]�h�j��  j  K	ubK
j	  )��}�(h�K$j  ]�h�j��  j  K
ubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubKj	  )��}�(h�K$j  ]�h�j��  j  KubK j	  )��}�(h�K$j  ]�h�j��  j  K ubK!j	  )��}�(h�K$j  ]�h�j��  j  K!ubK"j	  )��}�(h�K$j  ]�h�j��  j  K"ubK#j	  )��}�(h�K$j  ]�h�j��  j  K#ubK$j	  )��}�(h�K$j  ]�h�j��  j  K$ubK%j	  )��}�(h�K$j  ]�h�j��  j  K%ubK&j	  )��}�(h�K$j  ]�h�j��  j  K&ubK'j	  )��}�(h�K$j  ]�h�j��  j  K'ubK(j	  )��}�(h�K$j  ]�h�j��  j  K(ubK)j	  )��}�(h�K$j  ]�h�j��  j  K)ubK*j	  )��}�(h�K$j  ]�h�j��  j  K*ubK+j	  )��}�(h�K$j  ]�h�j��  j  K+ubK,j	  )��}�(h�K$j  ]�h�j��  j  K,ubK-j	  )��}�(h�K$j  ]�h�j��  j  K-ubK.j	  )��}�(h�K$j  ]�h�j��  j  K.ubK/j	  )��}�(h�K$j  ]�h�j��  j  K/ubK0j	  )��}�(h�K$j  ]�h�j��  j  K0ubK1j	  )��}�(h�K$j  ]�h�j��  j  K1ubK2j	  )��}�(h�K$j  ]�h�j��  j  K2ubK3j	  )��}�(h�K$j  ]�h�j��  j  K3ubK4j	  )��}�(h�K$j  ]�h�j��  j  K4ubK5j	  )��}�(h�K$j  ]�h�j��  j  K5ubK6j	  )��}�(h�K$j  ]�h�j��  j  K6ubK7j	  )��}�(h�K$j  ]�h�j��  j  K7ubK8j	  )��}�(h�K$j  ]�h�j��  j  K8ubK9j	  )��}�(h�K$j  ]�h�j��  j  K9ubK:j	  )��}�(h�K$j  ]�h�j��  j  K:ubK;j	  )��}�(h�K$j  ]�h�j��  j  K;ubK<j	  )��}�(h�K$j  ]�h�j��  j  K<ubK=j	  )��}�(h�K$j  ]�h�j��  j  K=ubK>j	  )��}�(h�K$j  ]�h�j��  j  K>ubK?j	  )��}�(h�K$j  ]�Kah�j��  j  K?ubK@j	  )��}�(h�K$j  ]�h�j��  j  K@ubKAj	  )��}�(h�K$j  ]�h�j��  j  KAubKBj	  )��}�(h�K$j  ]�h�j��  j  KBubKCj	  )��}�(h�K$j  ]�h�j��  j  KCubuK%}�(K j	  )��}�(h�K%j  ]�h�j��  j  K ubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubK	j	  )��}�(h�K%j  ]�h�j��  j  K	ubK
j	  )��}�(h�K%j  ]�h�j��  j  K
ubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubKj	  )��}�(h�K%j  ]�h�j��  j  KubK j	  )��}�(h�K%j  ]�h�j��  j  K ubK!j	  )��}�(h�K%j  ]�h�j��  j  K!ubK"j	  )��}�(h�K%j  ]�h�j��  j  K"ubK#j	  )��}�(h�K%j  ]�h�j��  j  K#ubK$j	  )��}�(h�K%j  ]�h�j��  j  K$ubK%j	  )��}�(h�K%j  ]�h�j��  j  K%ubK&j	  )��}�(h�K%j  ]�h�j��  j  K&ubK'j	  )��}�(h�K%j  ]�h�j��  j  K'ubK(j	  )��}�(h�K%j  ]�h�j��  j  K(ubK)j	  )��}�(h�K%j  ]�h�j��  j  K)ubK*j	  )��}�(h�K%j  ]�h�j��  j  K*ubK+j	  )��}�(h�K%j  ]�h�j��  j  K+ubK,j	  )��}�(h�K%j  ]�h�j��  j  K,ubK-j	  )��}�(h�K%j  ]�h�j��  j  K-ubK.j	  )��}�(h�K%j  ]�h�j��  j  K.ubK/j	  )��}�(h�K%j  ]�h�j��  j  K/ubK0j	  )��}�(h�K%j  ]�h�j��  j  K0ubK1j	  )��}�(h�K%j  ]�h�j��  j  K1ubK2j	  )��}�(h�K%j  ]�h�j��  j  K2ubK3j	  )��}�(h�K%j  ]�h�j��  j  K3ubK4j	  )��}�(h�K%j  ]�h�j��  j  K4ubK5j	  )��}�(h�K%j  ]�h�j��  j  K5ubK6j	  )��}�(h�K%j  ]�h�j��  j  K6ubK7j	  )��}�(h�K%j  ]�h�j��  j  K7ubK8j	  )��}�(h�K%j  ]�h�j��  j  K8ubK9j	  )��}�(h�K%j  ]�h�j��  j  K9ubK:j	  )��}�(h�K%j  ]�h�j��  j  K:ubK;j	  )��}�(h�K%j  ]�h�j��  j  K;ubK<j	  )��}�(h�K%j  ]�h�j��  j  K<ubK=j	  )��}�(h�K%j  ]�h�j��  j  K=ubK>j	  )��}�(h�K%j  ]�h�j��  j  K>ubK?j	  )��}�(h�K%j  ]�h�j��  j  K?ubK@j	  )��}�(h�K%j  ]�h�j��  j  K@ubKAj	  )��}�(h�K%j  ]�h�j��  j  KAubKBj	  )��}�(h�K%j  ]�h�j��  j  KBubKCj	  )��}�(h�K%j  ]�h�j��  j  KCubuK&}�(K j	  )��}�(h�K&j  ]�h�j��  j  K ubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubK	j	  )��}�(h�K&j  ]�h�j��  j  K	ubK
j	  )��}�(h�K&j  ]�h�j��  j  K
ubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubKj	  )��}�(h�K&j  ]�h�j��  j  KubK j	  )��}�(h�K&j  ]�h�j��  j  K ubK!j	  )��}�(h�K&j  ]�h�j��  j  K!ubK"j	  )��}�(h�K&j  ]�h�j��  j  K"ubK#j	  )��}�(h�K&j  ]�h�j��  j  K#ubK$j	  )��}�(h�K&j  ]�h�j��  j  K$ubK%j	  )��}�(h�K&j  ]�h�j��  j  K%ubK&j	  )��}�(h�K&j  ]�h�j��  j  K&ubK'j	  )��}�(h�K&j  ]�h�j��  j  K'ubK(j	  )��}�(h�K&j  ]�h�j��  j  K(ubK)j	  )��}�(h�K&j  ]�h�j��  j  K)ubK*j	  )��}�(h�K&j  ]�h�j��  j  K*ubK+j	  )��}�(h�K&j  ]�h�j��  j  K+ubK,j	  )��}�(h�K&j  ]�h�j��  j  K,ubK-j	  )��}�(h�K&j  ]�h�j��  j  K-ubK.j	  )��}�(h�K&j  ]�h�j��  j  K.ubK/j	  )��}�(h�K&j  ]�h�j��  j  K/ubK0j	  )��}�(h�K&j  ]�h�j��  j  K0ubK1j	  )��}�(h�K&j  ]�h�j��  j  K1ubK2j	  )��}�(h�K&j  ]�h�j��  j  K2ubK3j	  )��}�(h�K&j  ]�h�j��  j  K3ubK4j	  )��}�(h�K&j  ]�h�j��  j  K4ubK5j	  )��}�(h�K&j  ]�h�j��  j  K5ubK6j	  )��}�(h�K&j  ]�h�j��  j  K6ubK7j	  )��}�(h�K&j  ]�h�j��  j  K7ubK8j	  )��}�(h�K&j  ]�h�j��  j  K8ubK9j	  )��}�(h�K&j  ]�h�j��  j  K9ubK:j	  )��}�(h�K&j  ]�h�j��  j  K:ubK;j	  )��}�(h�K&j  ]�h�j��  j  K;ubK<j	  )��}�(h�K&j  ]�h�j��  j  K<ubK=j	  )��}�(h�K&j  ]�h�j��  j  K=ubK>j	  )��}�(h�K&j  ]�h�j��  j  K>ubK?j	  )��}�(h�K&j  ]�h�j��  j  K?ubK@j	  )��}�(h�K&j  ]�h�j��  j  K@ubKAj	  )��}�(h�K&j  ]�h�j��  j  KAubKBj	  )��}�(h�K&j  ]�h�j��  j  KBubKCj	  )��}�(h�K&j  ]�h�j��  j  KCubuK'}�(K j	  )��}�(h�K'j  ]�h�j��  j  K ubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubK	j	  )��}�(h�K'j  ]�h�j��  j  K	ubK
j	  )��}�(h�K'j  ]�h�j��  j  K
ubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubKj	  )��}�(h�K'j  ]�h�j��  j  KubK j	  )��}�(h�K'j  ]�h�j��  j  K ubK!j	  )��}�(h�K'j  ]�h�j��  j  K!ubK"j	  )��}�(h�K'j  ]�h�j��  j  K"ubK#j	  )��}�(h�K'j  ]�h�j��  j  K#ubK$j	  )��}�(h�K'j  ]�h�j��  j  K$ubK%j	  )��}�(h�K'j  ]�h�j��  j  K%ubK&j	  )��}�(h�K'j  ]�h�j��  j  K&ubK'j	  )��}�(h�K'j  ]�h�j��  j  K'ubK(j	  )��}�(h�K'j  ]�h�j��  j  K(ubK)j	  )��}�(h�K'j  ]�h�j��  j  K)ubK*j	  )��}�(h�K'j  ]�h�j��  j  K*ubK+j	  )��}�(h�K'j  ]�h�j��  j  K+ubK,j	  )��}�(h�K'j  ]�h�j��  j  K,ubK-j	  )��}�(h�K'j  ]�h�j��  j  K-ubK.j	  )��}�(h�K'j  ]�h�j��  j  K.ubK/j	  )��}�(h�K'j  ]�h�j��  j  K/ubK0j	  )��}�(h�K'j  ]�h�j��  j  K0ubK1j	  )��}�(h�K'j  ]�h�j��  j  K1ubK2j	  )��}�(h�K'j  ]�h�j��  j  K2ubK3j	  )��}�(h�K'j  ]�h�j��  j  K3ubK4j	  )��}�(h�K'j  ]�h�j��  j  K4ubK5j	  )��}�(h�K'j  ]�h�j��  j  K5ubK6j	  )��}�(h�K'j  ]�h�j��  j  K6ubK7j	  )��}�(h�K'j  ]�h�j��  j  K7ubK8j	  )��}�(h�K'j  ]�h�j��  j  K8ubK9j	  )��}�(h�K'j  ]�h�j��  j  K9ubK:j	  )��}�(h�K'j  ]�h�j��  j  K:ubK;j	  )��}�(h�K'j  ]�h�j��  j  K;ubK<j	  )��}�(h�K'j  ]�h�j��  j  K<ubK=j	  )��}�(h�K'j  ]�h�j��  j  K=ubK>j	  )��}�(h�K'j  ]�h�j��  j  K>ubK?j	  )��}�(h�K'j  ]�h�j��  j  K?ubK@j	  )��}�(h�K'j  ]�h�j��  j  K@ubKAj	  )��}�(h�K'j  ]�h�j��  j  KAubKBj	  )��}�(h�K'j  ]�h�j��  j  KBubKCj	  )��}�(h�K'j  ]�h�j��  j  KCubuK(}�(K j	  )��}�(h�K(j  ]�h�j��  j  K ubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubK	j	  )��}�(h�K(j  ]�h�j��  j  K	ubK
j	  )��}�(h�K(j  ]�h�j��  j  K
ubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubKj	  )��}�(h�K(j  ]�h�j��  j  KubK j	  )��}�(h�K(j  ]�h�j��  j  K ubK!j	  )��}�(h�K(j  ]�h�j��  j  K!ubK"j	  )��}�(h�K(j  ]�h�j��  j  K"ubK#j	  )��}�(h�K(j  ]�h�j��  j  K#ubK$j	  )��}�(h�K(j  ]�h�j��  j  K$ubK%j	  )��}�(h�K(j  ]�h�j��  j  K%ubK&j	  )��}�(h�K(j  ]�h�j��  j  K&ubK'j	  )��}�(h�K(j  ]�h�j��  j  K'ubK(j	  )��}�(h�K(j  ]�h�j��  j  K(ubK)j	  )��}�(h�K(j  ]�h�j��  j  K)ubK*j	  )��}�(h�K(j  ]�h�j��  j  K*ubK+j	  )��}�(h�K(j  ]�h�j��  j  K+ubK,j	  )��}�(h�K(j  ]�h�j��  j  K,ubK-j	  )��}�(h�K(j  ]�h�j��  j  K-ubK.j	  )��}�(h�K(j  ]�h�j��  j  K.ubK/j	  )��}�(h�K(j  ]�h�j��  j  K/ubK0j	  )��}�(h�K(j  ]�h�j��  j  K0ubK1j	  )��}�(h�K(j  ]�h�j��  j  K1ubK2j	  )��}�(h�K(j  ]�h�j��  j  K2ubK3j	  )��}�(h�K(j  ]�h�j��  j  K3ubK4j	  )��}�(h�K(j  ]�h�j��  j  K4ubK5j	  )��}�(h�K(j  ]�h�j��  j  K5ubK6j	  )��}�(h�K(j  ]�h�j��  j  K6ubK7j	  )��}�(h�K(j  ]�h�j��  j  K7ubK8j	  )��}�(h�K(j  ]�h�j��  j  K8ubK9j	  )��}�(h�K(j  ]�h�j��  j  K9ubK:j	  )��}�(h�K(j  ]�h�j��  j  K:ubK;j	  )��}�(h�K(j  ]�h�j��  j  K;ubK<j	  )��}�(h�K(j  ]�h�j��  j  K<ubK=j	  )��}�(h�K(j  ]�h�j��  j  K=ubK>j	  )��}�(h�K(j  ]�h�j��  j  K>ubK?j	  )��}�(h�K(j  ]�h�j��  j  K?ubK@j	  )��}�(h�K(j  ]�h�j��  j  K@ubKAj	  )��}�(h�K(j  ]�h�j��  j  KAubKBj	  )��}�(h�K(j  ]�h�j��  j  KBubKCj	  )��}�(h�K(j  ]�h�j��  j  KCubuK)}�(K j	  )��}�(h�K)j  ]�h�j��  j  K ubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubK	j	  )��}�(h�K)j  ]�h�j��  j  K	ubK
j	  )��}�(h�K)j  ]�h�j��  j  K
ubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubKj	  )��}�(h�K)j  ]�h�j��  j  KubK j	  )��}�(h�K)j  ]�h�j��  j  K ubK!j	  )��}�(h�K)j  ]�h�j��  j  K!ubK"j	  )��}�(h�K)j  ]�h�j��  j  K"ubK#j	  )��}�(h�K)j  ]�h�j��  j  K#ubK$j	  )��}�(h�K)j  ]�h�j��  j  K$ubK%j	  )��}�(h�K)j  ]�h�j��  j  K%ubK&j	  )��}�(h�K)j  ]�h�j��  j  K&ubK'j	  )��}�(h�K)j  ]�h�j��  j  K'ubK(j	  )��}�(h�K)j  ]�h�j��  j  K(ubK)j	  )��}�(h�K)j  ]�h�j��  j  K)ubK*j	  )��}�(h�K)j  ]�h�j��  j  K*ubK+j	  )��}�(h�K)j  ]�h�j��  j  K+ubK,j	  )��}�(h�K)j  ]�h�j��  j  K,ubK-j	  )��}�(h�K)j  ]�h�j��  j  K-ubK.j	  )��}�(h�K)j  ]�h�j��  j  K.ubK/j	  )��}�(h�K)j  ]�h�j��  j  K/ubK0j	  )��}�(h�K)j  ]�h�j��  j  K0ubK1j	  )��}�(h�K)j  ]�h�j��  j  K1ubK2j	  )��}�(h�K)j  ]�h�j��  j  K2ubK3j	  )��}�(h�K)j  ]�h�j��  j  K3ubK4j	  )��}�(h�K)j  ]�h�j��  j  K4ubK5j	  )��}�(h�K)j  ]�h�j��  j  K5ubK6j	  )��}�(h�K)j  ]�h�j��  j  K6ubK7j	  )��}�(h�K)j  ]�h�j��  j  K7ubK8j	  )��}�(h�K)j  ]�h�j��  j  K8ubK9j	  )��}�(h�K)j  ]�h�j��  j  K9ubK:j	  )��}�(h�K)j  ]�h�j��  j  K:ubK;j	  )��}�(h�K)j  ]�h�j��  j  K;ubK<j	  )��}�(h�K)j  ]�h�j��  j  K<ubK=j	  )��}�(h�K)j  ]�h�j��  j  K=ubK>j	  )��}�(h�K)j  ]�h�j��  j  K>ubK?j	  )��}�(h�K)j  ]�h�j��  j  K?ubK@j	  )��}�(h�K)j  ]�h�j��  j  K@ubKAj	  )��}�(h�K)j  ]�h�j��  j  KAubKBj	  )��}�(h�K)j  ]�h�j��  j  KBubKCj	  )��}�(h�K)j  ]�h�j��  j  KCubuK*}�(K j	  )��}�(h�K*j  ]�h�j��  j  K ubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubK	j	  )��}�(h�K*j  ]�h�j��  j  K	ubK
j	  )��}�(h�K*j  ]�h�j��  j  K
ubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubKj	  )��}�(h�K*j  ]�h�j��  j  KubK j	  )��}�(h�K*j  ]�h�j��  j  K ubK!j	  )��}�(h�K*j  ]�h�j��  j  K!ubK"j	  )��}�(h�K*j  ]�h�j��  j  K"ubK#j	  )��}�(h�K*j  ]�h�j��  j  K#ubK$j	  )��}�(h�K*j  ]�h�j��  j  K$ubK%j	  )��}�(h�K*j  ]�h�j��  j  K%ubK&j	  )��}�(h�K*j  ]�h�j��  j  K&ubK'j	  )��}�(h�K*j  ]�h�j��  j  K'ubK(j	  )��}�(h�K*j  ]�h�j��  j  K(ubK)j	  )��}�(h�K*j  ]�h�j��  j  K)ubK*j	  )��}�(h�K*j  ]�h�j��  j  K*ubK+j	  )��}�(h�K*j  ]�h�j��  j  K+ubK,j	  )��}�(h�K*j  ]�h�j��  j  K,ubK-j	  )��}�(h�K*j  ]�h�j��  j  K-ubK.j	  )��}�(h�K*j  ]�h�j��  j  K.ubK/j	  )��}�(h�K*j  ]�h�j��  j  K/ubK0j	  )��}�(h�K*j  ]�h�j��  j  K0ubK1j	  )��}�(h�K*j  ]�h�j��  j  K1ubK2j	  )��}�(h�K*j  ]�h�j��  j  K2ubK3j	  )��}�(h�K*j  ]�h�j��  j  K3ubK4j	  )��}�(h�K*j  ]�h�j��  j  K4ubK5j	  )��}�(h�K*j  ]�h�j��  j  K5ubK6j	  )��}�(h�K*j  ]�h�j��  j  K6ubK7j	  )��}�(h�K*j  ]�h�j��  j  K7ubK8j	  )��}�(h�K*j  ]�h�j��  j  K8ubK9j	  )��}�(h�K*j  ]�h�j��  j  K9ubK:j	  )��}�(h�K*j  ]�h�j��  j  K:ubK;j	  )��}�(h�K*j  ]�h�j��  j  K;ubK<j	  )��}�(h�K*j  ]�h�j��  j  K<ubK=j	  )��}�(h�K*j  ]�h�j��  j  K=ubK>j	  )��}�(h�K*j  ]�h�j��  j  K>ubK?j	  )��}�(h�K*j  ]�h�j��  j  K?ubK@j	  )��}�(h�K*j  ]�h�j��  j  K@ubKAj	  )��}�(h�K*j  ]�h�j��  j  KAubKBj	  )��}�(h�K*j  ]�h�j��  j  KBubKCj	  )��}�(h�K*j  ]�h�j��  j  KCubuK+}�(K j	  )��}�(h�K+j  ]�h�j��  j  K ubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubK	j	  )��}�(h�K+j  ]�h�j��  j  K	ubK
j	  )��}�(h�K+j  ]�h�j��  j  K
ubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubKj	  )��}�(h�K+j  ]�h�j��  j  KubK j	  )��}�(h�K+j  ]�h�j��  j  K ubK!j	  )��}�(h�K+j  ]�h�j��  j  K!ubK"j	  )��}�(h�K+j  ]�h�j��  j  K"ubK#j	  )��}�(h�K+j  ]�h�j��  j  K#ubK$j	  )��}�(h�K+j  ]�h�j��  j  K$ubK%j	  )��}�(h�K+j  ]�h�j��  j  K%ubK&j	  )��}�(h�K+j  ]�h�j��  j  K&ubK'j	  )��}�(h�K+j  ]�h�j��  j  K'ubK(j	  )��}�(h�K+j  ]�h�j��  j  K(ubK)j	  )��}�(h�K+j  ]�h�j��  j  K)ubK*j	  )��}�(h�K+j  ]�h�j��  j  K*ubK+j	  )��}�(h�K+j  ]�h�j��  j  K+ubK,j	  )��}�(h�K+j  ]�h�j��  j  K,ubK-j	  )��}�(h�K+j  ]�h�j��  j  K-ubK.j	  )��}�(h�K+j  ]�h�j��  j  K.ubK/j	  )��}�(h�K+j  ]�h�j��  j  K/ubK0j	  )��}�(h�K+j  ]�h�j��  j  K0ubK1j	  )��}�(h�K+j  ]�h�j��  j  K1ubK2j	  )��}�(h�K+j  ]�h�j��  j  K2ubK3j	  )��}�(h�K+j  ]�h�j��  j  K3ubK4j	  )��}�(h�K+j  ]�h�j��  j  K4ubK5j	  )��}�(h�K+j  ]�h�j��  j  K5ubK6j	  )��}�(h�K+j  ]�h�j��  j  K6ubK7j	  )��}�(h�K+j  ]�h�j��  j  K7ubK8j	  )��}�(h�K+j  ]�h�j��  j  K8ubK9j	  )��}�(h�K+j  ]�h�j��  j  K9ubK:j	  )��}�(h�K+j  ]�h�j��  j  K:ubK;j	  )��}�(h�K+j  ]�h�j��  j  K;ubK<j	  )��}�(h�K+j  ]�h�j��  j  K<ubK=j	  )��}�(h�K+j  ]�h�j��  j  K=ubK>j	  )��}�(h�K+j  ]�h�j��  j  K>ubK?j	  )��}�(h�K+j  ]�h�j��  j  K?ubK@j	  )��}�(h�K+j  ]�h�j��  j  K@ubKAj	  )��}�(h�K+j  ]�h�j��  j  KAubKBj	  )��}�(h�K+j  ]�h�j��  j  KBubKCj	  )��}�(h�K+j  ]�h�j��  j  KCubuK,}�(K j	  )��}�(h�K,j  ]�h�j��  j  K ubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubK	j	  )��}�(h�K,j  ]�h�j��  j  K	ubK
j	  )��}�(h�K,j  ]�h�j��  j  K
ubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubKj	  )��}�(h�K,j  ]�h�j��  j  KubK j	  )��}�(h�K,j  ]�h�j��  j  K ubK!j	  )��}�(h�K,j  ]�h�j��  j  K!ubK"j	  )��}�(h�K,j  ]�h�j��  j  K"ubK#j	  )��}�(h�K,j  ]�h�j��  j  K#ubK$j	  )��}�(h�K,j  ]�h�j��  j  K$ubK%j	  )��}�(h�K,j  ]�h�j��  j  K%ubK&j	  )��}�(h�K,j  ]�h�j��  j  K&ubK'j	  )��}�(h�K,j  ]�h�j��  j  K'ubK(j	  )��}�(h�K,j  ]�h�j��  j  K(ubK)j	  )��}�(h�K,j  ]�h�j��  j  K)ubK*j	  )��}�(h�K,j  ]�h�j��  j  K*ubK+j	  )��}�(h�K,j  ]�h�j��  j  K+ubK,j	  )��}�(h�K,j  ]�h�j��  j  K,ubK-j	  )��}�(h�K,j  ]�h�j��  j  K-ubK.j	  )��}�(h�K,j  ]�h�j��  j  K.ubK/j	  )��}�(h�K,j  ]�h�j��  j  K/ubK0j	  )��}�(h�K,j  ]�h�j��  j  K0ubK1j	  )��}�(h�K,j  ]�h�j��  j  K1ubK2j	  )��}�(h�K,j  ]�h�j��  j  K2ubK3j	  )��}�(h�K,j  ]�h�j��  j  K3ubK4j	  )��}�(h�K,j  ]�h�j��  j  K4ubK5j	  )��}�(h�K,j  ]�h�j��  j  K5ubK6j	  )��}�(h�K,j  ]�h�j��  j  K6ubK7j	  )��}�(h�K,j  ]�h�j��  j  K7ubK8j	  )��}�(h�K,j  ]�h�j��  j  K8ubK9j	  )��}�(h�K,j  ]�h�j��  j  K9ubK:j	  )��}�(h�K,j  ]�h�j��  j  K:ubK;j	  )��}�(h�K,j  ]�h�j��  j  K;ubK<j	  )��}�(h�K,j  ]�h�j��  j  K<ubK=j	  )��}�(h�K,j  ]�h�j��  j  K=ubK>j	  )��}�(h�K,j  ]�h�j��  j  K>ubK?j	  )��}�(h�K,j  ]�h�j��  j  K?ubK@j	  )��}�(h�K,j  ]�h�j��  j  K@ubKAj	  )��}�(h�K,j  ]�h�j��  j  KAubKBj	  )��}�(h�K,j  ]�h�j��  j  KBubKCj	  )��}�(h�K,j  ]�h�j��  j  KCubuK-}�(K j	  )��}�(h�K-j  ]�h�j��  j  K ubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubK	j	  )��}�(h�K-j  ]�h�j��  j  K	ubK
j	  )��}�(h�K-j  ]�h�j��  j  K
ubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubKj	  )��}�(h�K-j  ]�h�j��  j  KubK j	  )��}�(h�K-j  ]�h�j��  j  K ubK!j	  )��}�(h�K-j  ]�h�j��  j  K!ubK"j	  )��}�(h�K-j  ]�h�j��  j  K"ubK#j	  )��}�(h�K-j  ]�h�j��  j  K#ubK$j	  )��}�(h�K-j  ]�h�j��  j  K$ubK%j	  )��}�(h�K-j  ]�h�j��  j  K%ubK&j	  )��}�(h�K-j  ]�h�j��  j  K&ubK'j	  )��}�(h�K-j  ]�h�j��  j  K'ubK(j	  )��}�(h�K-j  ]�h�j��  j  K(ubK)j	  )��}�(h�K-j  ]�h�j��  j  K)ubK*j	  )��}�(h�K-j  ]�h�j��  j  K*ubK+j	  )��}�(h�K-j  ]�h�j��  j  K+ubK,j	  )��}�(h�K-j  ]�h�j��  j  K,ubK-j	  )��}�(h�K-j  ]�h�j��  j  K-ubK.j	  )��}�(h�K-j  ]�h�j��  j  K.ubK/j	  )��}�(h�K-j  ]�h�j��  j  K/ubK0j	  )��}�(h�K-j  ]�h�j��  j  K0ubK1j	  )��}�(h�K-j  ]�h�j��  j  K1ubK2j	  )��}�(h�K-j  ]�h�j��  j  K2ubK3j	  )��}�(h�K-j  ]�h�j��  j  K3ubK4j	  )��}�(h�K-j  ]�h�j��  j  K4ubK5j	  )��}�(h�K-j  ]�h�j��  j  K5ubK6j	  )��}�(h�K-j  ]�h�j��  j  K6ubK7j	  )��}�(h�K-j  ]�h�j��  j  K7ubK8j	  )��}�(h�K-j  ]�h�j��  j  K8ubK9j	  )��}�(h�K-j  ]�h�j��  j  K9ubK:j	  )��}�(h�K-j  ]�h�j��  j  K:ubK;j	  )��}�(h�K-j  ]�h�j��  j  K;ubK<j	  )��}�(h�K-j  ]�h�j��  j  K<ubK=j	  )��}�(h�K-j  ]�h�j��  j  K=ubK>j	  )��}�(h�K-j  ]�h�j��  j  K>ubK?j	  )��}�(h�K-j  ]�h�j��  j  K?ubK@j	  )��}�(h�K-j  ]�h�j��  j  K@ubKAj	  )��}�(h�K-j  ]�h�j��  j  KAubKBj	  )��}�(h�K-j  ]�h�j��  j  KBubKCj	  )��}�(h�K-j  ]�h�j��  j  KCubuK.}�(K j	  )��}�(h�K.j  ]�h�j��  j  K ubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubK	j	  )��}�(h�K.j  ]�h�j��  j  K	ubK
j	  )��}�(h�K.j  ]�h�j��  j  K
ubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubKj	  )��}�(h�K.j  ]�h�j��  j  KubK j	  )��}�(h�K.j  ]�h�j��  j  K ubK!j	  )��}�(h�K.j  ]�h�j��  j  K!ubK"j	  )��}�(h�K.j  ]�h�j��  j  K"ubK#j	  )��}�(h�K.j  ]�h�j��  j  K#ubK$j	  )��}�(h�K.j  ]�h�j��  j  K$ubK%j	  )��}�(h�K.j  ]�h�j��  j  K%ubK&j	  )��}�(h�K.j  ]�h�j��  j  K&ubK'j	  )��}�(h�K.j  ]�h�j��  j  K'ubK(j	  )��}�(h�K.j  ]�h�j��  j  K(ubK)j	  )��}�(h�K.j  ]�h�j��  j  K)ubK*j	  )��}�(h�K.j  ]�h�j��  j  K*ubK+j	  )��}�(h�K.j  ]�h�j��  j  K+ubK,j	  )��}�(h�K.j  ]�h�j��  j  K,ubK-j	  )��}�(h�K.j  ]�h�j��  j  K-ubK.j	  )��}�(h�K.j  ]�h�j��  j  K.ubK/j	  )��}�(h�K.j  ]�h�j��  j  K/ubK0j	  )��}�(h�K.j  ]�h�j��  j  K0ubK1j	  )��}�(h�K.j  ]�h�j��  j  K1ubK2j	  )��}�(h�K.j  ]�h�j��  j  K2ubK3j	  )��}�(h�K.j  ]�h�j��  j  K3ubK4j	  )��}�(h�K.j  ]�h�j��  j  K4ubK5j	  )��}�(h�K.j  ]�h�j��  j  K5ubK6j	  )��}�(h�K.j  ]�h�j��  j  K6ubK7j	  )��}�(h�K.j  ]�h�j��  j  K7ubK8j	  )��}�(h�K.j  ]�h�j��  j  K8ubK9j	  )��}�(h�K.j  ]�h�j��  j  K9ubK:j	  )��}�(h�K.j  ]�h�j��  j  K:ubK;j	  )��}�(h�K.j  ]�h�j��  j  K;ubK<j	  )��}�(h�K.j  ]�h�j��  j  K<ubK=j	  )��}�(h�K.j  ]�h�j��  j  K=ubK>j	  )��}�(h�K.j  ]�h�j��  j  K>ubK?j	  )��}�(h�K.j  ]�h�j��  j  K?ubK@j	  )��}�(h�K.j  ]�h�j��  j  K@ubKAj	  )��}�(h�K.j  ]�h�j��  j  KAubKBj	  )��}�(h�K.j  ]�h�j��  j  KBubKCj	  )��}�(h�K.j  ]�h�j��  j  KCubuK/}�(K j	  )��}�(h�K/j  ]�h�j��  j  K ubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubK	j	  )��}�(h�K/j  ]�h�j��  j  K	ubK
j	  )��}�(h�K/j  ]�h�j��  j  K
ubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubKj	  )��}�(h�K/j  ]�h�j��  j  KubK j	  )��}�(h�K/j  ]�h�j��  j  K ubK!j	  )��}�(h�K/j  ]�h�j��  j  K!ubK"j	  )��}�(h�K/j  ]�h�j��  j  K"ubK#j	  )��}�(h�K/j  ]�h�j��  j  K#ubK$j	  )��}�(h�K/j  ]�h�j��  j  K$ubK%j	  )��}�(h�K/j  ]�h�j��  j  K%ubK&j	  )��}�(h�K/j  ]�h�j��  j  K&ubK'j	  )��}�(h�K/j  ]�h�j��  j  K'ubK(j	  )��}�(h�K/j  ]�h�j��  j  K(ubK)j	  )��}�(h�K/j  ]�h�j��  j  K)ubK*j	  )��}�(h�K/j  ]�h�j��  j  K*ubK+j	  )��}�(h�K/j  ]�h�j��  j  K+ubK,j	  )��}�(h�K/j  ]�h�j��  j  K,ubK-j	  )��}�(h�K/j  ]�h�j��  j  K-ubK.j	  )��}�(h�K/j  ]�h�j��  j  K.ubK/j	  )��}�(h�K/j  ]�h�j��  j  K/ubK0j	  )��}�(h�K/j  ]�h�j��  j  K0ubK1j	  )��}�(h�K/j  ]�h�j��  j  K1ubK2j	  )��}�(h�K/j  ]�h�j��  j  K2ubK3j	  )��}�(h�K/j  ]�h�j��  j  K3ubK4j	  )��}�(h�K/j  ]�h�j��  j  K4ubK5j	  )��}�(h�K/j  ]�h�j��  j  K5ubK6j	  )��}�(h�K/j  ]�h�j��  j  K6ubK7j	  )��}�(h�K/j  ]�h�j��  j  K7ubK8j	  )��}�(h�K/j  ]�h�j��  j  K8ubK9j	  )��}�(h�K/j  ]�h�j��  j  K9ubK:j	  )��}�(h�K/j  ]�h�j��  j  K:ubK;j	  )��}�(h�K/j  ]�h�j��  j  K;ubK<j	  )��}�(h�K/j  ]�h�j��  j  K<ubK=j	  )��}�(h�K/j  ]�h�j��  j  K=ubK>j	  )��}�(h�K/j  ]�h�j��  j  K>ubK?j	  )��}�(h�K/j  ]�h�j��  j  K?ubK@j	  )��}�(h�K/j  ]�h�j��  j  K@ubKAj	  )��}�(h�K/j  ]�h�j��  j  KAubKBj	  )��}�(h�K/j  ]�h�j��  j  KBubKCj	  )��}�(h�K/j  ]�h�j��  j  KCubuK0}�(K j	  )��}�(h�K0j  ]�h�j��  j  K ubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubK	j	  )��}�(h�K0j  ]�h�j��  j  K	ubK
j	  )��}�(h�K0j  ]�h�j��  j  K
ubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubKj	  )��}�(h�K0j  ]�h�j��  j  KubK j	  )��}�(h�K0j  ]�h�j��  j  K ubK!j	  )��}�(h�K0j  ]�h�j��  j  K!ubK"j	  )��}�(h�K0j  ]�h�j��  j  K"ubK#j	  )��}�(h�K0j  ]�h�j��  j  K#ubK$j	  )��}�(h�K0j  ]�h�j��  j  K$ubK%j	  )��}�(h�K0j  ]�h�j��  j  K%ubK&j	  )��}�(h�K0j  ]�h�j��  j  K&ubK'j	  )��}�(h�K0j  ]�h�j��  j  K'ubK(j	  )��}�(h�K0j  ]�h�j��  j  K(ubK)j	  )��}�(h�K0j  ]�h�j��  j  K)ubK*j	  )��}�(h�K0j  ]�h�j��  j  K*ubK+j	  )��}�(h�K0j  ]�h�j��  j  K+ubK,j	  )��}�(h�K0j  ]�h�j��  j  K,ubK-j	  )��}�(h�K0j  ]�h�j��  j  K-ubK.j	  )��}�(h�K0j  ]�h�j��  j  K.ubK/j	  )��}�(h�K0j  ]�h�j��  j  K/ubK0j	  )��}�(h�K0j  ]�h�j��  j  K0ubK1j	  )��}�(h�K0j  ]�h�j��  j  K1ubK2j	  )��}�(h�K0j  ]�h�j��  j  K2ubK3j	  )��}�(h�K0j  ]�h�j��  j  K3ubK4j	  )��}�(h�K0j  ]�h�j��  j  K4ubK5j	  )��}�(h�K0j  ]�h�j��  j  K5ubK6j	  )��}�(h�K0j  ]�h�j��  j  K6ubK7j	  )��}�(h�K0j  ]�h�j��  j  K7ubK8j	  )��}�(h�K0j  ]�h�j��  j  K8ubK9j	  )��}�(h�K0j  ]�h�j��  j  K9ubK:j	  )��}�(h�K0j  ]�h�j��  j  K:ubK;j	  )��}�(h�K0j  ]�h�j��  j  K;ubK<j	  )��}�(h�K0j  ]�h�j��  j  K<ubK=j	  )��}�(h�K0j  ]�h�j��  j  K=ubK>j	  )��}�(h�K0j  ]�h�j��  j  K>ubK?j	  )��}�(h�K0j  ]�h�j��  j  K?ubK@j	  )��}�(h�K0j  ]�h�j��  j  K@ubKAj	  )��}�(h�K0j  ]�h�j��  j  KAubKBj	  )��}�(h�K0j  ]�h�j��  j  KBubKCj	  )��}�(h�K0j  ]�h�j��  j  KCubuK1}�(K j	  )��}�(h�K1j  ]�h�j��  j  K ubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubK	j	  )��}�(h�K1j  ]�h�j��  j  K	ubK
j	  )��}�(h�K1j  ]�h�j��  j  K
ubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubKj	  )��}�(h�K1j  ]�h�j��  j  KubK j	  )��}�(h�K1j  ]�h�j��  j  K ubK!j	  )��}�(h�K1j  ]�h�j��  j  K!ubK"j	  )��}�(h�K1j  ]�h�j��  j  K"ubK#j	  )��}�(h�K1j  ]�h�j��  j  K#ubK$j	  )��}�(h�K1j  ]�h�j��  j  K$ubK%j	  )��}�(h�K1j  ]�h�j��  j  K%ubK&j	  )��}�(h�K1j  ]�h�j��  j  K&ubK'j	  )��}�(h�K1j  ]�h�j��  j  K'ubK(j	  )��}�(h�K1j  ]�h�j��  j  K(ubK)j	  )��}�(h�K1j  ]�h�j��  j  K)ubK*j	  )��}�(h�K1j  ]�h�j��  j  K*ubK+j	  )��}�(h�K1j  ]�h�j��  j  K+ubK,j	  )��}�(h�K1j  ]�h�j��  j  K,ubK-j	  )��}�(h�K1j  ]�h�j��  j  K-ubK.j	  )��}�(h�K1j  ]�h�j��  j  K.ubK/j	  )��}�(h�K1j  ]�h�j��  j  K/ubK0j	  )��}�(h�K1j  ]�h�j��  j  K0ubK1j	  )��}�(h�K1j  ]�h�j��  j  K1ubK2j	  )��}�(h�K1j  ]�h�j��  j  K2ubK3j	  )��}�(h�K1j  ]�h�j��  j  K3ubK4j	  )��}�(h�K1j  ]�h�j��  j  K4ubK5j	  )��}�(h�K1j  ]�h�j��  j  K5ubK6j	  )��}�(h�K1j  ]�h�j��  j  K6ubK7j	  )��}�(h�K1j  ]�h�j��  j  K7ubK8j	  )��}�(h�K1j  ]�h�j��  j  K8ubK9j	  )��}�(h�K1j  ]�h�j��  j  K9ubK:j	  )��}�(h�K1j  ]�h�j��  j  K:ubK;j	  )��}�(h�K1j  ]�h�j��  j  K;ubK<j	  )��}�(h�K1j  ]�h�j��  j  K<ubK=j	  )��}�(h�K1j  ]�h�j��  j  K=ubK>j	  )��}�(h�K1j  ]�h�j��  j  K>ubK?j	  )��}�(h�K1j  ]�h�j��  j  K?ubK@j	  )��}�(h�K1j  ]�h�j��  j  K@ubKAj	  )��}�(h�K1j  ]�h�j��  j  KAubKBj	  )��}�(h�K1j  ]�h�j��  j  KBubKCj	  )��}�(h�K1j  ]�h�j��  j  KCubuK2}�(K j	  )��}�(h�K2j  ]�h�j��  j  K ubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubK	j	  )��}�(h�K2j  ]�h�j��  j  K	ubK
j	  )��}�(h�K2j  ]�h�j��  j  K
ubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubKj	  )��}�(h�K2j  ]�h�j��  j  KubK j	  )��}�(h�K2j  ]�h�j��  j  K ubK!j	  )��}�(h�K2j  ]�h�j��  j  K!ubK"j	  )��}�(h�K2j  ]�h�j��  j  K"ubK#j	  )��}�(h�K2j  ]�h�j��  j  K#ubK$j	  )��}�(h�K2j  ]�h�j��  j  K$ubK%j	  )��}�(h�K2j  ]�h�j��  j  K%ubK&j	  )��}�(h�K2j  ]�h�j��  j  K&ubK'j	  )��}�(h�K2j  ]�h�j��  j  K'ubK(j	  )��}�(h�K2j  ]�h�j��  j  K(ubK)j	  )��}�(h�K2j  ]�h�j��  j  K)ubK*j	  )��}�(h�K2j  ]�h�j��  j  K*ubK+j	  )��}�(h�K2j  ]�h�j��  j  K+ubK,j	  )��}�(h�K2j  ]�h�j��  j  K,ubK-j	  )��}�(h�K2j  ]�h�j��  j  K-ubK.j	  )��}�(h�K2j  ]�h�j��  j  K.ubK/j	  )��}�(h�K2j  ]�h�j��  j  K/ubK0j	  )��}�(h�K2j  ]�h�j��  j  K0ubK1j	  )��}�(h�K2j  ]�h�j��  j  K1ubK2j	  )��}�(h�K2j  ]�h�j��  j  K2ubK3j	  )��}�(h�K2j  ]�h�j��  j  K3ubK4j	  )��}�(h�K2j  ]�h�j��  j  K4ubK5j	  )��}�(h�K2j  ]�h�j��  j  K5ubK6j	  )��}�(h�K2j  ]�h�j��  j  K6ubK7j	  )��}�(h�K2j  ]�h�j��  j  K7ubK8j	  )��}�(h�K2j  ]�h�j��  j  K8ubK9j	  )��}�(h�K2j  ]�h�j��  j  K9ubK:j	  )��}�(h�K2j  ]�h�j��  j  K:ubK;j	  )��}�(h�K2j  ]�h�j��  j  K;ubK<j	  )��}�(h�K2j  ]�h�j��  j  K<ubK=j	  )��}�(h�K2j  ]�h�j��  j  K=ubK>j	  )��}�(h�K2j  ]�h�j��  j  K>ubK?j	  )��}�(h�K2j  ]�h�j��  j  K?ubK@j	  )��}�(h�K2j  ]�h�j��  j  K@ubKAj	  )��}�(h�K2j  ]�h�j��  j  KAubKBj	  )��}�(h�K2j  ]�h�j��  j  KBubKCj	  )��}�(h�K2j  ]�h�j��  j  KCubuK3}�(K j	  )��}�(h�K3j  ]�h�j��  j  K ubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubK	j	  )��}�(h�K3j  ]�h�j��  j  K	ubK
j	  )��}�(h�K3j  ]�h�j��  j  K
ubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubKj	  )��}�(h�K3j  ]�h�j��  j  KubK j	  )��}�(h�K3j  ]�h�j��  j  K ubK!j	  )��}�(h�K3j  ]�h�j��  j  K!ubK"j	  )��}�(h�K3j  ]�h�j��  j  K"ubK#j	  )��}�(h�K3j  ]�h�j��  j  K#ubK$j	  )��}�(h�K3j  ]�h�j��  j  K$ubK%j	  )��}�(h�K3j  ]�h�j��  j  K%ubK&j	  )��}�(h�K3j  ]�h�j��  j  K&ubK'j	  )��}�(h�K3j  ]�h�j��  j  K'ubK(j	  )��}�(h�K3j  ]�h�j��  j  K(ubK)j	  )��}�(h�K3j  ]�h�j��  j  K)ubK*j	  )��}�(h�K3j  ]�h�j��  j  K*ubK+j	  )��}�(h�K3j  ]�h�j��  j  K+ubK,j	  )��}�(h�K3j  ]�h�j��  j  K,ubK-j	  )��}�(h�K3j  ]�h�j��  j  K-ubK.j	  )��}�(h�K3j  ]�h�j��  j  K.ubK/j	  )��}�(h�K3j  ]�h�j��  j  K/ubK0j	  )��}�(h�K3j  ]�h�j��  j  K0ubK1j	  )��}�(h�K3j  ]�h�j��  j  K1ubK2j	  )��}�(h�K3j  ]�h�j��  j  K2ubK3j	  )��}�(h�K3j  ]�h�j��  j  K3ubK4j	  )��}�(h�K3j  ]�h�j��  j  K4ubK5j	  )��}�(h�K3j  ]�h�j��  j  K5ubK6j	  )��}�(h�K3j  ]�h�j��  j  K6ubK7j	  )��}�(h�K3j  ]�h�j��  j  K7ubK8j	  )��}�(h�K3j  ]�h�j��  j  K8ubK9j	  )��}�(h�K3j  ]�h�j��  j  K9ubK:j	  )��}�(h�K3j  ]�h�j��  j  K:ubK;j	  )��}�(h�K3j  ]�h�j��  j  K;ubK<j	  )��}�(h�K3j  ]�h�j��  j  K<ubK=j	  )��}�(h�K3j  ]�h�j��  j  K=ubK>j	  )��}�(h�K3j  ]�h�j��  j  K>ubK?j	  )��}�(h�K3j  ]�h�j��  j  K?ubK@j	  )��}�(h�K3j  ]�h�j��  j  K@ubKAj	  )��}�(h�K3j  ]�h�j��  j  KAubKBj	  )��}�(h�K3j  ]�h�j��  j  KBubKCj	  )��}�(h�K3j  ]�h�j��  j  KCubuK4}�(K j	  )��}�(h�K4j  ]�h�j��  j  K ubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubK	j	  )��}�(h�K4j  ]�h�j��  j  K	ubK
j	  )��}�(h�K4j  ]�h�j��  j  K
ubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubKj	  )��}�(h�K4j  ]�h�j��  j  KubK j	  )��}�(h�K4j  ]�h�j��  j  K ubK!j	  )��}�(h�K4j  ]�h�j��  j  K!ubK"j	  )��}�(h�K4j  ]�h�j��  j  K"ubK#j	  )��}�(h�K4j  ]�h�j��  j  K#ubK$j	  )��}�(h�K4j  ]�h�j��  j  K$ubK%j	  )��}�(h�K4j  ]�h�j��  j  K%ubK&j	  )��}�(h�K4j  ]�h�j��  j  K&ubK'j	  )��}�(h�K4j  ]�h�j��  j  K'ubK(j	  )��}�(h�K4j  ]�h�j��  j  K(ubK)j	  )��}�(h�K4j  ]�h�j��  j  K)ubK*j	  )��}�(h�K4j  ]�h�j��  j  K*ubK+j	  )��}�(h�K4j  ]�h�j��  j  K+ubK,j	  )��}�(h�K4j  ]�h�j��  j  K,ubK-j	  )��}�(h�K4j  ]�h�j��  j  K-ubK.j	  )��}�(h�K4j  ]�h�j��  j  K.ubK/j	  )��}�(h�K4j  ]�h�j��  j  K/ubK0j	  )��}�(h�K4j  ]�h�j��  j  K0ubK1j	  )��}�(h�K4j  ]�h�j��  j  K1ubK2j	  )��}�(h�K4j  ]�h�j��  j  K2ubK3j	  )��}�(h�K4j  ]�h�j��  j  K3ubK4j	  )��}�(h�K4j  ]�h�j��  j  K4ubK5j	  )��}�(h�K4j  ]�h�j��  j  K5ubK6j	  )��}�(h�K4j  ]�h�j��  j  K6ubK7j	  )��}�(h�K4j  ]�h�j��  j  K7ubK8j	  )��}�(h�K4j  ]�h�j��  j  K8ubK9j	  )��}�(h�K4j  ]�h�j��  j  K9ubK:j	  )��}�(h�K4j  ]�h�j��  j  K:ubK;j	  )��}�(h�K4j  ]�h�j��  j  K;ubK<j	  )��}�(h�K4j  ]�h�j��  j  K<ubK=j	  )��}�(h�K4j  ]�h�j��  j  K=ubK>j	  )��}�(h�K4j  ]�h�j��  j  K>ubK?j	  )��}�(h�K4j  ]�h�j��  j  K?ubK@j	  )��}�(h�K4j  ]�h�j��  j  K@ubKAj	  )��}�(h�K4j  ]�h�j��  j  KAubKBj	  )��}�(h�K4j  ]�h�j��  j  KBubKCj	  )��}�(h�K4j  ]�h�j��  j  KCubuK5}�(K j	  )��}�(h�K5j  ]�h�j��  j  K ubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubK	j	  )��}�(h�K5j  ]�h�j��  j  K	ubK
j	  )��}�(h�K5j  ]�h�j��  j  K
ubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubKj	  )��}�(h�K5j  ]�h�j��  j  KubK j	  )��}�(h�K5j  ]�h�j��  j  K ubK!j	  )��}�(h�K5j  ]�h�j��  j  K!ubK"j	  )��}�(h�K5j  ]�h�j��  j  K"ubK#j	  )��}�(h�K5j  ]�h�j��  j  K#ubK$j	  )��}�(h�K5j  ]�h�j��  j  K$ubK%j	  )��}�(h�K5j  ]�h�j��  j  K%ubK&j	  )��}�(h�K5j  ]�h�j��  j  K&ubK'j	  )��}�(h�K5j  ]�h�j��  j  K'ubK(j	  )��}�(h�K5j  ]�h�j��  j  K(ubK)j	  )��}�(h�K5j  ]�h�j��  j  K)ubK*j	  )��}�(h�K5j  ]�h�j��  j  K*ubK+j	  )��}�(h�K5j  ]�h�j��  j  K+ubK,j	  )��}�(h�K5j  ]�h�j��  j  K,ubK-j	  )��}�(h�K5j  ]�h�j��  j  K-ubK.j	  )��}�(h�K5j  ]�h�j��  j  K.ubK/j	  )��}�(h�K5j  ]�h�j��  j  K/ubK0j	  )��}�(h�K5j  ]�h�j��  j  K0ubK1j	  )��}�(h�K5j  ]�h�j��  j  K1ubK2j	  )��}�(h�K5j  ]�h�j��  j  K2ubK3j	  )��}�(h�K5j  ]�h�j��  j  K3ubK4j	  )��}�(h�K5j  ]�h�j��  j  K4ubK5j	  )��}�(h�K5j  ]�h�j��  j  K5ubK6j	  )��}�(h�K5j  ]�h�j��  j  K6ubK7j	  )��}�(h�K5j  ]�h�j��  j  K7ubK8j	  )��}�(h�K5j  ]�h�j��  j  K8ubK9j	  )��}�(h�K5j  ]�h�j��  j  K9ubK:j	  )��}�(h�K5j  ]�h�j��  j  K:ubK;j	  )��}�(h�K5j  ]�h�j��  j  K;ubK<j	  )��}�(h�K5j  ]�h�j��  j  K<ubK=j	  )��}�(h�K5j  ]�Kah�j��  j  K=ubK>j	  )��}�(h�K5j  ]�h�j��  j  K>ubK?j	  )��}�(h�K5j  ]�h�j��  j  K?ubK@j	  )��}�(h�K5j  ]�h�j��  j  K@ubKAj	  )��}�(h�K5j  ]�h�j��  j  KAubKBj	  )��}�(h�K5j  ]�h�j��  j  KBubKCj	  )��}�(h�K5j  ]�h�j��  j  KCubuK6}�(K j	  )��}�(h�K6j  ]�h�j��  j  K ubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubK	j	  )��}�(h�K6j  ]�h�j��  j  K	ubK
j	  )��}�(h�K6j  ]�h�j��  j  K
ubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubKj	  )��}�(h�K6j  ]�h�j��  j  KubK j	  )��}�(h�K6j  ]�h�j��  j  K ubK!j	  )��}�(h�K6j  ]�h�j��  j  K!ubK"j	  )��}�(h�K6j  ]�h�j��  j  K"ubK#j	  )��}�(h�K6j  ]�h�j��  j  K#ubK$j	  )��}�(h�K6j  ]�h�j��  j  K$ubK%j	  )��}�(h�K6j  ]�h�j��  j  K%ubK&j	  )��}�(h�K6j  ]�h�j��  j  K&ubK'j	  )��}�(h�K6j  ]�h�j��  j  K'ubK(j	  )��}�(h�K6j  ]�h�j��  j  K(ubK)j	  )��}�(h�K6j  ]�h�j��  j  K)ubK*j	  )��}�(h�K6j  ]�h�j��  j  K*ubK+j	  )��}�(h�K6j  ]�h�j��  j  K+ubK,j	  )��}�(h�K6j  ]�h�j��  j  K,ubK-j	  )��}�(h�K6j  ]�h�j��  j  K-ubK.j	  )��}�(h�K6j  ]�h�j��  j  K.ubK/j	  )��}�(h�K6j  ]�h�j��  j  K/ubK0j	  )��}�(h�K6j  ]�h�j��  j  K0ubK1j	  )��}�(h�K6j  ]�h�j��  j  K1ubK2j	  )��}�(h�K6j  ]�h�j��  j  K2ubK3j	  )��}�(h�K6j  ]�h�j��  j  K3ubK4j	  )��}�(h�K6j  ]�h�j��  j  K4ubK5j	  )��}�(h�K6j  ]�h�j��  j  K5ubK6j	  )��}�(h�K6j  ]�h�j��  j  K6ubK7j	  )��}�(h�K6j  ]�h�j��  j  K7ubK8j	  )��}�(h�K6j  ]�h�j��  j  K8ubK9j	  )��}�(h�K6j  ]�h�j��  j  K9ubK:j	  )��}�(h�K6j  ]�h�j��  j  K:ubK;j	  )��}�(h�K6j  ]�h�j��  j  K;ubK<j	  )��}�(h�K6j  ]�h�j��  j  K<ubK=j	  )��}�(h�K6j  ]�h�j��  j  K=ubK>j	  )��}�(h�K6j  ]�h�j��  j  K>ubK?j	  )��}�(h�K6j  ]�h�j��  j  K?ubK@j	  )��}�(h�K6j  ]�h�j��  j  K@ubKAj	  )��}�(h�K6j  ]�h�j��  j  KAubKBj	  )��}�(h�K6j  ]�h�j��  j  KBubKCj	  )��}�(h�K6j  ]�h�j��  j  KCubuK7}�(K j	  )��}�(h�K7j  ]�h�j��  j  K ubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubK	j	  )��}�(h�K7j  ]�h�j��  j  K	ubK
j	  )��}�(h�K7j  ]�h�j��  j  K
ubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubKj	  )��}�(h�K7j  ]�h�j��  j  KubK j	  )��}�(h�K7j  ]�h�j��  j  K ubK!j	  )��}�(h�K7j  ]�h�j��  j  K!ubK"j	  )��}�(h�K7j  ]�h�j��  j  K"ubK#j	  )��}�(h�K7j  ]�h�j��  j  K#ubK$j	  )��}�(h�K7j  ]�h�j��  j  K$ubK%j	  )��}�(h�K7j  ]�h�j��  j  K%ubK&j	  )��}�(h�K7j  ]�h�j��  j  K&ubK'j	  )��}�(h�K7j  ]�h�j��  j  K'ubK(j	  )��}�(h�K7j  ]�h�j��  j  K(ubK)j	  )��}�(h�K7j  ]�h�j��  j  K)ubK*j	  )��}�(h�K7j  ]�h�j��  j  K*ubK+j	  )��}�(h�K7j  ]�h�j��  j  K+ubK,j	  )��}�(h�K7j  ]�h�j��  j  K,ubK-j	  )��}�(h�K7j  ]�h�j��  j  K-ubK.j	  )��}�(h�K7j  ]�h�j��  j  K.ubK/j	  )��}�(h�K7j  ]�h�j��  j  K/ubK0j	  )��}�(h�K7j  ]�h�j��  j  K0ubK1j	  )��}�(h�K7j  ]�h�j��  j  K1ubK2j	  )��}�(h�K7j  ]�h�j��  j  K2ubK3j	  )��}�(h�K7j  ]�h�j��  j  K3ubK4j	  )��}�(h�K7j  ]�h�j��  j  K4ubK5j	  )��}�(h�K7j  ]�h�j��  j  K5ubK6j	  )��}�(h�K7j  ]�h�j��  j  K6ubK7j	  )��}�(h�K7j  ]�h�j��  j  K7ubK8j	  )��}�(h�K7j  ]�h�j��  j  K8ubK9j	  )��}�(h�K7j  ]�h�j��  j  K9ubK:j	  )��}�(h�K7j  ]�h�j��  j  K:ubK;j	  )��}�(h�K7j  ]�h�j��  j  K;ubK<j	  )��}�(h�K7j  ]�h�j��  j  K<ubK=j	  )��}�(h�K7j  ]�Kah�j��  j  K=ubK>j	  )��}�(h�K7j  ]�h�j��  j  K>ubK?j	  )��}�(h�K7j  ]�h�j��  j  K?ubK@j	  )��}�(h�K7j  ]�Kah�j��  j  K@ubKAj	  )��}�(h�K7j  ]�h�j��  j  KAubKBj	  )��}�(h�K7j  ]�h�j��  j  KBubKCj	  )��}�(h�K7j  ]�h�j��  j  KCubuK8}�(K j	  )��}�(h�K8j  ]�h�j��  j  K ubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubK	j	  )��}�(h�K8j  ]�h�j��  j  K	ubK
j	  )��}�(h�K8j  ]�h�j��  j  K
ubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubKj	  )��}�(h�K8j  ]�h�j��  j  KubK j	  )��}�(h�K8j  ]�h�j��  j  K ubK!j	  )��}�(h�K8j  ]�h�j��  j  K!ubK"j	  )��}�(h�K8j  ]�h�j��  j  K"ubK#j	  )��}�(h�K8j  ]�h�j��  j  K#ubK$j	  )��}�(h�K8j  ]�h�j��  j  K$ubK%j	  )��}�(h�K8j  ]�h�j��  j  K%ubK&j	  )��}�(h�K8j  ]�h�j��  j  K&ubK'j	  )��}�(h�K8j  ]�h�j��  j  K'ubK(j	  )��}�(h�K8j  ]�h�j��  j  K(ubK)j	  )��}�(h�K8j  ]�h�j��  j  K)ubK*j	  )��}�(h�K8j  ]�h�j��  j  K*ubK+j	  )��}�(h�K8j  ]�h�j��  j  K+ubK,j	  )��}�(h�K8j  ]�h�j��  j  K,ubK-j	  )��}�(h�K8j  ]�h�j��  j  K-ubK.j	  )��}�(h�K8j  ]�h�j��  j  K.ubK/j	  )��}�(h�K8j  ]�h�j��  j  K/ubK0j	  )��}�(h�K8j  ]�h�j��  j  K0ubK1j	  )��}�(h�K8j  ]�h�j��  j  K1ubK2j	  )��}�(h�K8j  ]�h�j��  j  K2ubK3j	  )��}�(h�K8j  ]�h�j��  j  K3ubK4j	  )��}�(h�K8j  ]�h�j��  j  K4ubK5j	  )��}�(h�K8j  ]�h�j��  j  K5ubK6j	  )��}�(h�K8j  ]�h�j��  j  K6ubK7j	  )��}�(h�K8j  ]�h�j��  j  K7ubK8j	  )��}�(h�K8j  ]�h�j��  j  K8ubK9j	  )��}�(h�K8j  ]�h�j��  j  K9ubK:j	  )��}�(h�K8j  ]�h�j��  j  K:ubK;j	  )��}�(h�K8j  ]�h�j��  j  K;ubK<j	  )��}�(h�K8j  ]�h�j��  j  K<ubK=j	  )��}�(h�K8j  ]�h�j��  j  K=ubK>j	  )��}�(h�K8j  ]�h�j��  j  K>ubK?j	  )��}�(h�K8j  ]�h�j��  j  K?ubK@j	  )��}�(h�K8j  ]�h�j��  j  K@ubKAj	  )��}�(h�K8j  ]�h�j��  j  KAubKBj	  )��}�(h�K8j  ]�h�j��  j  KBubKCj	  )��}�(h�K8j  ]�h�j��  j  KCubuK9}�(K j	  )��}�(h�K9j  ]�h�j��  j  K ubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubK	j	  )��}�(h�K9j  ]�h�j��  j  K	ubK
j	  )��}�(h�K9j  ]�h�j��  j  K
ubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubKj	  )��}�(h�K9j  ]�h�j��  j  KubK j	  )��}�(h�K9j  ]�h�j��  j  K ubK!j	  )��}�(h�K9j  ]�h�j��  j  K!ubK"j	  )��}�(h�K9j  ]�h�j��  j  K"ubK#j	  )��}�(h�K9j  ]�h�j��  j  K#ubK$j	  )��}�(h�K9j  ]�h�j��  j  K$ubK%j	  )��}�(h�K9j  ]�h�j��  j  K%ubK&j	  )��}�(h�K9j  ]�h�j��  j  K&ubK'j	  )��}�(h�K9j  ]�h�j��  j  K'ubK(j	  )��}�(h�K9j  ]�h�j��  j  K(ubK)j	  )��}�(h�K9j  ]�h�j��  j  K)ubK*j	  )��}�(h�K9j  ]�h�j��  j  K*ubK+j	  )��}�(h�K9j  ]�h�j��  j  K+ubK,j	  )��}�(h�K9j  ]�h�j��  j  K,ubK-j	  )��}�(h�K9j  ]�h�j��  j  K-ubK.j	  )��}�(h�K9j  ]�h�j��  j  K.ubK/j	  )��}�(h�K9j  ]�h�j��  j  K/ubK0j	  )��}�(h�K9j  ]�h�j��  j  K0ubK1j	  )��}�(h�K9j  ]�h�j��  j  K1ubK2j	  )��}�(h�K9j  ]�h�j��  j  K2ubK3j	  )��}�(h�K9j  ]�h�j��  j  K3ubK4j	  )��}�(h�K9j  ]�h�j��  j  K4ubK5j	  )��}�(h�K9j  ]�h�j��  j  K5ubK6j	  )��}�(h�K9j  ]�h�j��  j  K6ubK7j	  )��}�(h�K9j  ]�h�j��  j  K7ubK8j	  )��}�(h�K9j  ]�h�j��  j  K8ubK9j	  )��}�(h�K9j  ]�h�j��  j  K9ubK:j	  )��}�(h�K9j  ]�h�j��  j  K:ubK;j	  )��}�(h�K9j  ]�h�j��  j  K;ubK<j	  )��}�(h�K9j  ]�h�j��  j  K<ubK=j	  )��}�(h�K9j  ]�h�j��  j  K=ubK>j	  )��}�(h�K9j  ]�h�j��  j  K>ubK?j	  )��}�(h�K9j  ]�h�j��  j  K?ubK@j	  )��}�(h�K9j  ]�h�j��  j  K@ubKAj	  )��}�(h�K9j  ]�h�j��  j  KAubKBj	  )��}�(h�K9j  ]�h�j��  j  KBubKCj	  )��}�(h�K9j  ]�h�j��  j  KCubuK:}�(K j	  )��}�(h�K:j  ]�h�j��  j  K ubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubK	j	  )��}�(h�K:j  ]�h�j��  j  K	ubK
j	  )��}�(h�K:j  ]�h�j��  j  K
ubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  �      KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubKj	  )��}�(h�K:j  ]�h�j��  j  KubK j	  )��}�(h�K:j  ]�h�j��  j  K ubK!j	  )��}�(h�K:j  ]�h�j��  j  K!ubK"j	  )��}�(h�K:j  ]�h�j��  j  K"ubK#j	  )��}�(h�K:j  ]�h�j��  j  K#ubK$j	  )��}�(h�K:j  ]�h�j��  j  K$ubK%j	  )��}�(h�K:j  ]�h�j��  j  K%ubK&j	  )��}�(h�K:j  ]�h�j��  j  K&ubK'j	  )��}�(h�K:j  ]�h�j��  j  K'ubK(j	  )��}�(h�K:j  ]�h�j��  j  K(ubK)j	  )��}�(h�K:j  ]�h�j��  j  K)ubK*j	  )��}�(h�K:j  ]�h�j��  j  K*ubK+j	  )��}�(h�K:j  ]�h�j��  j  K+ubK,j	  )��}�(h�K:j  ]�h�j��  j  K,ubK-j	  )��}�(h�K:j  ]�h�j��  j  K-ubK.j	  )��}�(h�K:j  ]�h�j��  j  K.ubK/j	  )��}�(h�K:j  ]�h�j��  j  K/ubK0j	  )��}�(h�K:j  ]�h�j��  j  K0ubK1j	  )��}�(h�K:j  ]�h�j��  j  K1ubK2j	  )��}�(h�K:j  ]�h�j��  j  K2ubK3j	  )��}�(h�K:j  ]�h�j��  j  K3ubK4j	  )��}�(h�K:j  ]�h�j��  j  K4ubK5j	  )��}�(h�K:j  ]�h�j��  j  K5ubK6j	  )��}�(h�K:j  ]�h�j��  j  K6ubK7j	  )��}�(h�K:j  ]�h�j��  j  K7ubK8j	  )��}�(h�K:j  ]�h�j��  j  K8ubK9j	  )��}�(h�K:j  ]�h�j��  j  K9ubK:j	  )��}�(h�K:j  ]�h�j��  j  K:ubK;j	  )��}�(h�K:j  ]�h�j��  j  K;ubK<j	  )��}�(h�K:j  ]�h�j��  j  K<ubK=j	  )��}�(h�K:j  ]�h�j��  j  K=ubK>j	  )��}�(h�K:j  ]�h�j��  j  K>ubK?j	  )��}�(h�K:j  ]�h�j��  j  K?ubK@j	  )��}�(h�K:j  ]�h�j��  j  K@ubKAj	  )��}�(h�K:j  ]�h�j��  j  KAubKBj	  )��}�(h�K:j  ]�h�j��  j  KBubKCj	  )��}�(h�K:j  ]�h�j��  j  KCubuK;}�(K j	  )��}�(h�K;j  ]�h�j��  j  K ubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�Kah�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubK	j	  )��}�(h�K;j  ]�h�j��  j  K	ubK
j	  )��}�(h�K;j  ]�h�j��  j  K
ubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubKj	  )��}�(h�K;j  ]�h�j��  j  KubK j	  )��}�(h�K;j  ]�h�j��  j  K ubK!j	  )��}�(h�K;j  ]�h�j��  j  K!ubK"j	  )��}�(h�K;j  ]�h�j��  j  K"ubK#j	  )��}�(h�K;j  ]�h�j��  j  K#ubK$j	  )��}�(h�K;j  ]�h�j��  j  K$ubK%j	  )��}�(h�K;j  ]�h�j��  j  K%ubK&j	  )��}�(h�K;j  ]�h�j��  j  K&ubK'j	  )��}�(h�K;j  ]�h�j��  j  K'ubK(j	  )��}�(h�K;j  ]�h�j��  j  K(ubK)j	  )��}�(h�K;j  ]�h�j��  j  K)ubK*j	  )��}�(h�K;j  ]�h�j��  j  K*ubK+j	  )��}�(h�K;j  ]�h�j��  j  K+ubK,j	  )��}�(h�K;j  ]�h�j��  j  K,ubK-j	  )��}�(h�K;j  ]�h�j��  j  K-ubK.j	  )��}�(h�K;j  ]�h�j��  j  K.ubK/j	  )��}�(h�K;j  ]�h�j��  j  K/ubK0j	  )��}�(h�K;j  ]�h�j��  j  K0ubK1j	  )��}�(h�K;j  ]�h�j��  j  K1ubK2j	  )��}�(h�K;j  ]�h�j��  j  K2ubK3j	  )��}�(h�K;j  ]�h�j��  j  K3ubK4j	  )��}�(h�K;j  ]�h�j��  j  K4ubK5j	  )��}�(h�K;j  ]�h�j��  j  K5ubK6j	  )��}�(h�K;j  ]�h�j��  j  K6ubK7j	  )��}�(h�K;j  ]�h�j��  j  K7ubK8j	  )��}�(h�K;j  ]�h�j��  j  K8ubK9j	  )��}�(h�K;j  ]�h�j��  j  K9ubK:j	  )��}�(h�K;j  ]�h�j��  j  K:ubK;j	  )��}�(h�K;j  ]�h�j��  j  K;ubK<j	  )��}�(h�K;j  ]�h�j��  j  K<ubK=j	  )��}�(h�K;j  ]�h�j��  j  K=ubK>j	  )��}�(h�K;j  ]�h�j��  j  K>ubK?j	  )��}�(h�K;j  ]�h�j��  j  K?ubK@j	  )��}�(h�K;j  ]�h�j��  j  K@ubKAj	  )��}�(h�K;j  ]�h�j��  j  KAubKBj	  )��}�(h�K;j  ]�h�j��  j  KBubKCj	  )��}�(h�K;j  ]�h�j��  j  KCubuK<}�(K j	  )��}�(h�K<j  ]�h�j��  j  K ubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubK	j	  )��}�(h�K<j  ]�h�j��  j  K	ubK
j	  )��}�(h�K<j  ]�h�j��  j  K
ubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�Kah�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubKj	  )��}�(h�K<j  ]�h�j��  j  KubK j	  )��}�(h�K<j  ]�h�j��  j  K ubK!j	  )��}�(h�K<j  ]�h�j��  j  K!ubK"j	  )��}�(h�K<j  ]�h�j��  j  K"ubK#j	  )��}�(h�K<j  ]�h�j��  j  K#ubK$j	  )��}�(h�K<j  ]�h�j��  j  K$ubK%j	  )��}�(h�K<j  ]�h�j��  j  K%ubK&j	  )��}�(h�K<j  ]�h�j��  j  K&ubK'j	  )��}�(h�K<j  ]�h�j��  j  K'ubK(j	  )��}�(h�K<j  ]�h�j��  j  K(ubK)j	  )��}�(h�K<j  ]�h�j��  j  K)ubK*j	  )��}�(h�K<j  ]�h�j��  j  K*ubK+j	  )��}�(h�K<j  ]�h�j��  j  K+ubK,j	  )��}�(h�K<j  ]�h�j��  j  K,ubK-j	  )��}�(h�K<j  ]�h�j��  j  K-ubK.j	  )��}�(h�K<j  ]�h�j��  j  K.ubK/j	  )��}�(h�K<j  ]�h�j��  j  K/ubK0j	  )��}�(h�K<j  ]�h�j��  j  K0ubK1j	  )��}�(h�K<j  ]�h�j��  j  K1ubK2j	  )��}�(h�K<j  ]�h�j��  j  K2ubK3j	  )��}�(h�K<j  ]�h�j��  j  K3ubK4j	  )��}�(h�K<j  ]�h�j��  j  K4ubK5j	  )��}�(h�K<j  ]�h�j��  j  K5ubK6j	  )��}�(h�K<j  ]�h�j��  j  K6ubK7j	  )��}�(h�K<j  ]�h�j��  j  K7ubK8j	  )��}�(h�K<j  ]�h�j��  j  K8ubK9j	  )��}�(h�K<j  ]�h�j��  j  K9ubK:j	  )��}�(h�K<j  ]�h�j��  j  K:ubK;j	  )��}�(h�K<j  ]�h�j��  j  K;ubK<j	  )��}�(h�K<j  ]�h�j��  j  K<ubK=j	  )��}�(h�K<j  ]�h�j��  j  K=ubK>j	  )��}�(h�K<j  ]�h�j��  j  K>ubK?j	  )��}�(h�K<j  ]�h�j��  j  K?ubK@j	  )��}�(h�K<j  ]�h�j��  j  K@ubKAj	  )��}�(h�K<j  ]�h�j��  j  KAubKBj	  )��}�(h�K<j  ]�h�j��  j  KBubKCj	  )��}�(h�K<j  ]�h�j��  j  KCubuK=}�(K j	  )��}�(h�K=j  ]�h�j��  j  K ubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�Kah�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubK	j	  )��}�(h�K=j  ]�h�j��  j  K	ubK
j	  )��}�(h�K=j  ]�h�j��  j  K
ubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�Kah�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�Kah�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubKj	  )��}�(h�K=j  ]�h�j��  j  KubK j	  )��}�(h�K=j  ]�h�j��  j  K ubK!j	  )��}�(h�K=j  ]�h�j��  j  K!ubK"j	  )��}�(h�K=j  ]�h�j��  j  K"ubK#j	  )��}�(h�K=j  ]�h�j��  j  K#ubK$j	  )��}�(h�K=j  ]�h�j��  j  K$ubK%j	  )��}�(h�K=j  ]�h�j��  j  K%ubK&j	  )��}�(h�K=j  ]�h�j��  j  K&ubK'j	  )��}�(h�K=j  ]�h�j��  j  K'ubK(j	  )��}�(h�K=j  ]�h�j��  j  K(ubK)j	  )��}�(h�K=j  ]�h�j��  j  K)ubK*j	  )��}�(h�K=j  ]�h�j��  j  K*ubK+j	  )��}�(h�K=j  ]�h�j��  j  K+ubK,j	  )��}�(h�K=j  ]�h�j��  j  K,ubK-j	  )��}�(h�K=j  ]�h�j��  j  K-ubK.j	  )��}�(h�K=j  ]�h�j��  j  K.ubK/j	  )��}�(h�K=j  ]�h�j��  j  K/ubK0j	  )��}�(h�K=j  ]�h�j��  j  K0ubK1j	  )��}�(h�K=j  ]�h�j��  j  K1ubK2j	  )��}�(h�K=j  ]�h�j��  j  K2ubK3j	  )��}�(h�K=j  ]�h�j��  j  K3ubK4j	  )��}�(h�K=j  ]�h�j��  j  K4ubK5j	  )��}�(h�K=j  ]�h�j��  j  K5ubK6j	  )��}�(h�K=j  ]�h�j��  j  K6ubK7j	  )��}�(h�K=j  ]�h�j��  j  K7ubK8j	  )��}�(h�K=j  ]�h�j��  j  K8ubK9j	  )��}�(h�K=j  ]�h�j��  j  K9ubK:j	  )��}�(h�K=j  ]�h�j��  j  K:ubK;j	  )��}�(h�K=j  ]�h�j��  j  K;ubK<j	  )��}�(h�K=j  ]�h�j��  j  K<ubK=j	  )��}�(h�K=j  ]�h�j��  j  K=ubK>j	  )��}�(h�K=j  ]�h�j��  j  K>ubK?j	  )��}�(h�K=j  ]�h�j��  j  K?ubK@j	  )��}�(h�K=j  ]�h�j��  j  K@ubKAj	  )��}�(h�K=j  ]�h�j��  j  KAubKBj	  )��}�(h�K=j  ]�h�j��  j  KBubKCj	  )��}�(h�K=j  ]�h�j��  j  KCubuK>}�(K j	  )��}�(h�K>j  ]�h�j��  j  K ubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�Kah�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubK	j	  )��}�(h�K>j  ]�h�j��  j  K	ubK
j	  )��}�(h�K>j  ]�h�j��  j  K
ubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�Kah�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubKj	  )��}�(h�K>j  ]�h�j��  j  KubK j	  )��}�(h�K>j  ]�h�j��  j  K ubK!j	  )��}�(h�K>j  ]�h�j��  j  K!ubK"j	  )��}�(h�K>j  ]�h�j��  j  K"ubK#j	  )��}�(h�K>j  ]�h�j��  j  K#ubK$j	  )��}�(h�K>j  ]�h�j��  j  K$ubK%j	  )��}�(h�K>j  ]�h�j��  j  K%ubK&j	  )��}�(h�K>j  ]�h�j��  j  K&ubK'j	  )��}�(h�K>j  ]�h�j��  j  K'ubK(j	  )��}�(h�K>j  ]�h�j��  j  K(ubK)j	  )��}�(h�K>j  ]�h�j��  j  K)ubK*j	  )��}�(h�K>j  ]�h�j��  j  K*ubK+j	  )��}�(h�K>j  ]�h�j��  j  K+ubK,j	  )��}�(h�K>j  ]�h�j��  j  K,ubK-j	  )��}�(h�K>j  ]�h�j��  j  K-ubK.j	  )��}�(h�K>j  ]�h�j��  j  K.ubK/j	  )��}�(h�K>j  ]�h�j��  j  K/ubK0j	  )��}�(h�K>j  ]�h�j��  j  K0ubK1j	  )��}�(h�K>j  ]�h�j��  j  K1ubK2j	  )��}�(h�K>j  ]�h�j��  j  K2ubK3j	  )��}�(h�K>j  ]�h�j��  j  K3ubK4j	  )��}�(h�K>j  ]�h�j��  j  K4ubK5j	  )��}�(h�K>j  ]�h�j��  j  K5ubK6j	  )��}�(h�K>j  ]�h�j��  j  K6ubK7j	  )��}�(h�K>j  ]�h�j��  j  K7ubK8j	  )��}�(h�K>j  ]�h�j��  j  K8ubK9j	  )��}�(h�K>j  ]�h�j��  j  K9ubK:j	  )��}�(h�K>j  ]�h�j��  j  K:ubK;j	  )��}�(h�K>j  ]�h�j��  j  K;ubK<j	  )��}�(h�K>j  ]�h�j��  j  K<ubK=j	  )��}�(h�K>j  ]�h�j��  j  K=ubK>j	  )��}�(h�K>j  ]�h�j��  j  K>ubK?j	  )��}�(h�K>j  ]�h�j��  j  K?ubK@j	  )��}�(h�K>j  ]�h�j��  j  K@ubKAj	  )��}�(h�K>j  ]�h�j��  j  KAubKBj	  )��}�(h�K>j  ]�h�j��  j  KBubKCj	  )��}�(h�K>j  ]�h�j��  j  KCubuK?}�(K j	  )��}�(h�K?j  ]�h�j��  j  K ubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubK	j	  )��}�(h�K?j  ]�h�j��  j  K	ubK
j	  )��}�(h�K?j  ]�h�j��  j  K
ubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�Kah�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubKj	  )��}�(h�K?j  ]�h�j��  j  KubK j	  )��}�(h�K?j  ]�h�j��  j  K ubK!j	  )��}�(h�K?j  ]�h�j��  j  K!ubK"j	  )��}�(h�K?j  ]�h�j��  j  K"ubK#j	  )��}�(h�K?j  ]�h�j��  j  K#ubK$j	  )��}�(h�K?j  ]�h�j��  j  K$ubK%j	  )��}�(h�K?j  ]�h�j��  j  K%ubK&j	  )��}�(h�K?j  ]�h�j��  j  K&ubK'j	  )��}�(h�K?j  ]�Kah�j��  j  K'ubK(j	  )��}�(h�K?j  ]�h�j��  j  K(ubK)j	  )��}�(h�K?j  ]�h�j��  j  K)ubK*j	  )��}�(h�K?j  ]�h�j��  j  K*ubK+j	  )��}�(h�K?j  ]�h�j��  j  K+ubK,j	  )��}�(h�K?j  ]�h�j��  j  K,ubK-j	  )��}�(h�K?j  ]�h�j��  j  K-ubK.j	  )��}�(h�K?j  ]�h�j��  j  K.ubK/j	  )��}�(h�K?j  ]�h�j��  j  K/ubK0j	  )��}�(h�K?j  ]�h�j��  j  K0ubK1j	  )��}�(h�K?j  ]�h�j��  j  K1ubK2j	  )��}�(h�K?j  ]�h�j��  j  K2ubK3j	  )��}�(h�K?j  ]�h�j��  j  K3ubK4j	  )��}�(h�K?j  ]�h�j��  j  K4ubK5j	  )��}�(h�K?j  ]�h�j��  j  K5ubK6j	  )��}�(h�K?j  ]�h�j��  j  K6ubK7j	  )��}�(h�K?j  ]�h�j��  j  K7ubK8j	  )��}�(h�K?j  ]�h�j��  j  K8ubK9j	  )��}�(h�K?j  ]�h�j��  j  K9ubK:j	  )��}�(h�K?j  ]�h�j��  j  K:ubK;j	  )��}�(h�K?j  ]�h�j��  j  K;ubK<j	  )��}�(h�K?j  ]�h�j��  j  K<ubK=j	  )��}�(h�K?j  ]�h�j��  j  K=ubK>j	  )��}�(h�K?j  ]�h�j��  j  K>ubK?j	  )��}�(h�K?j  ]�h�j��  j  K?ubK@j	  )��}�(h�K?j  ]�h�j��  j  K@ubKAj	  )��}�(h�K?j  ]�h�j��  j  KAubKBj	  )��}�(h�K?j  ]�h�j��  j  KBubKCj	  )��}�(h�K?j  ]�h�j��  j  KCubuK@}�(K j	  )��}�(h�K@j  ]�h�j��  j  K ubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubK	j	  )��}�(h�K@j  ]�h�j��  j  K	ubK
j	  )��}�(h�K@j  ]�h�j��  j  K
ubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubKj	  )��}�(h�K@j  ]�h�j��  j  KubK j	  )��}�(h�K@j  ]�h�j��  j  K ubK!j	  )��}�(h�K@j  ]�h�j��  j  K!ubK"j	  )��}�(h�K@j  ]�h�j��  j  K"ubK#j	  )��}�(h�K@j  ]�h�j��  j  K#ubK$j	  )��}�(h�K@j  ]�Kah�j��  j  K$ubK%j	  )��}�(h�K@j  ]�Kah�j��  j  K%ubK&j	  )��}�(h�K@j  ]�h�j��  j  K&ubK'j	  )��}�(h�K@j  ]�h�j��  j  K'ubK(j	  )��}�(h�K@j  ]�h�j��  j  K(ubK)j	  )��}�(h�K@j  ]�h�j��  j  K)ubK*j	  )��}�(h�K@j  ]�h�j��  j  K*ubK+j	  )��}�(h�K@j  ]�h�j��  j  K+ubK,j	  )��}�(h�K@j  ]�h�j��  j  K,ubK-j	  )��}�(h�K@j  ]�h�j��  j  K-ubK.j	  )��}�(h�K@j  ]�h�j��  j  K.ubK/j	  )��}�(h�K@j  ]�h�j��  j  K/ubK0j	  )��}�(h�K@j  ]�h�j��  j  K0ubK1j	  )��}�(h�K@j  ]�h�j��  j  K1ubK2j	  )��}�(h�K@j  ]�h�j��  j  K2ubK3j	  )��}�(h�K@j  ]�h�j��  j  K3ubK4j	  )��}�(h�K@j  ]�h�j��  j  K4ubK5j	  )��}�(h�K@j  ]�h�j��  j  K5ubK6j	  )��}�(h�K@j  ]�h�j��  j  K6ubK7j	  )��}�(h�K@j  ]�h�j��  j  K7ubK8j	  )��}�(h�K@j  ]�h�j��  j  K8ubK9j	  )��}�(h�K@j  ]�h�j��  j  K9ubK:j	  )��}�(h�K@j  ]�h�j��  j  K:ubK;j	  )��}�(h�K@j  ]�h�j��  j  K;ubK<j	  )��}�(h�K@j  ]�h�j��  j  K<ubK=j	  )��}�(h�K@j  ]�h�j��  j  K=ubK>j	  )��}�(h�K@j  ]�h�j��  j  K>ubK?j	  )��}�(h�K@j  ]�h�j��  j  K?ubK@j	  )��}�(h�K@j  ]�h�j��  j  K@ubKAj	  )��}�(h�K@j  ]�h�j��  j  KAubKBj	  )��}�(h�K@j  ]�h�j��  j  KBubKCj	  )��}�(h�K@j  ]�h�j��  j  KCubuKA}�(K j	  )��}�(h�KAj  ]�h�j��  j  K ubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubK	j	  )��}�(h�KAj  ]�h�j��  j  K	ubK
j	  )��}�(h�KAj  ]�h�j��  j  K
ubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubKj	  )��}�(h�KAj  ]�h�j��  j  KubK j	  )��}�(h�KAj  ]�h�j��  j  K ubK!j	  )��}�(h�KAj  ]�h�j��  j  K!ubK"j	  )��}�(h�KAj  ]�Kah�j��  j  K"ubK#j	  )��}�(h�KAj  ]�h�j��  j  K#ubK$j	  )��}�(h�KAj  ]�h�j��  j  K$ubK%j	  )��}�(h�KAj  ]�h�j��  j  K%ubK&j	  )��}�(h�KAj  ]�h�j��  j  K&ubK'j	  )��}�(h�KAj  ]�h�j��  j  K'ubK(j	  )��}�(h�KAj  ]�h�j��  j  K(ubK)j	  )��}�(h�KAj  ]�h�j��  j  K)ubK*j	  )��}�(h�KAj  ]�h�j��  j  K*ubK+j	  )��}�(h�KAj  ]�h�j��  j  K+ubK,j	  )��}�(h�KAj  ]�h�j��  j  K,ubK-j	  )��}�(h�KAj  ]�h�j��  j  K-ubK.j	  )��}�(h�KAj  ]�h�j��  j  K.ubK/j	  )��}�(h�KAj  ]�h�j��  j  K/ubK0j	  )��}�(h�KAj  ]�h�j��  j  K0ubK1j	  )��}�(h�KAj  ]�h�j��  j  K1ubK2j	  )��}�(h�KAj  ]�h�j��  j  K2ubK3j	  )��}�(h�KAj  ]�h�j��  j  K3ubK4j	  )��}�(h�KAj  ]�h�j��  j  K4ubK5j	  )��}�(h�KAj  ]�h�j��  j  K5ubK6j	  )��}�(h�KAj  ]�h�j��  j  K6ubK7j	  )��}�(h�KAj  ]�h�j��  j  K7ubK8j	  )��}�(h�KAj  ]�h�j��  j  K8ubK9j	  )��}�(h�KAj  ]�h�j��  j  K9ubK:j	  )��}�(h�KAj  ]�h�j��  j  K:ubK;j	  )��}�(h�KAj  ]�h�j��  j  K;ubK<j	  )��}�(h�KAj  ]�h�j��  j  K<ubK=j	  )��}�(h�KAj  ]�h�j��  j  K=ubK>j	  )��}�(h�KAj  ]�h�j��  j  K>ubK?j	  )��}�(h�KAj  ]�h�j��  j  K?ubK@j	  )��}�(h�KAj  ]�h�j��  j  K@ubKAj	  )��}�(h�KAj  ]�h�j��  j  KAubKBj	  )��}�(h�KAj  ]�h�j��  j  KBubKCj	  )��}�(h�KAj  ]�h�j��  j  KCubuKB}�(K j	  )��}�(h�KBj  ]�h�j��  j  K ubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubK	j	  )��}�(h�KBj  ]�h�j��  j  K	ubK
j	  )��}�(h�KBj  ]�h�j��  j  K
ubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubKj	  )��}�(h�KBj  ]�h�j��  j  KubK j	  )��}�(h�KBj  ]�h�j��  j  K ubK!j	  )��}�(h�KBj  ]�h�j��  j  K!ubK"j	  )��}�(h�KBj  ]�h�j��  j  K"ubK#j	  )��}�(h�KBj  ]�h�j��  j  K#ubK$j	  )��}�(h�KBj  ]�h�j��  j  K$ubK%j	  )��}�(h�KBj  ]�h�j��  j  K%ubK&j	  )��}�(h�KBj  ]�h�j��  j  K&ubK'j	  )��}�(h�KBj  ]�h�j��  j  K'ubK(j	  )��}�(h�KBj  ]�h�j��  j  K(ubK)j	  )��}�(h�KBj  ]�h�j��  j  K)ubK*j	  )��}�(h�KBj  ]�h�j��  j  K*ubK+j	  )��}�(h�KBj  ]�h�j��  j  K+ubK,j	  )��}�(h�KBj  ]�h�j��  j  K,ubK-j	  )��}�(h�KBj  ]�h�j��  j  K-ubK.j	  )��}�(h�KBj  ]�h�j��  j  K.ubK/j	  )��}�(h�KBj  ]�h�j��  j  K/ubK0j	  )��}�(h�KBj  ]�h�j��  j  K0ubK1j	  )��}�(h�KBj  ]�h�j��  j  K1ubK2j	  )��}�(h�KBj  ]�h�j��  j  K2ubK3j	  )��}�(h�KBj  ]�h�j��  j  K3ubK4j	  )��}�(h�KBj  ]�h�j��  j  K4ubK5j	  )��}�(h�KBj  ]�h�j��  j  K5ubK6j	  )��}�(h�KBj  ]�h�j��  j  K6ubK7j	  )��}�(h�KBj  ]�h�j��  j  K7ubK8j	  )��}�(h�KBj  ]�h�j��  j  K8ubK9j	  )��}�(h�KBj  ]�h�j��  j  K9ubK:j	  )��}�(h�KBj  ]�h�j��  j  K:ubK;j	  )��}�(h�KBj  ]�h�j��  j  K;ubK<j	  )��}�(h�KBj  ]�h�j��  j  K<ubK=j	  )��}�(h�KBj  ]�h�j��  j  K=ubK>j	  )��}�(h�KBj  ]�h�j��  j  K>ubK?j	  )��}�(h�KBj  ]�h�j��  j  K?ubK@j	  )��}�(h�KBj  ]�h�j��  j  K@ubKAj	  )��}�(h�KBj  ]�h�j��  j  KAubKBj	  )��}�(h�KBj  ]�h�j��  j  KBubKCj	  )��}�(h�KBj  ]�h�j��  j  KCubuKC}�(K j	  )��}�(h�KCj  ]�h�j��  j  K ubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubK	j	  )��}�(h�KCj  ]�h�j��  j  K	ubK
j	  )��}�(h�KCj  ]�h�j��  j  K
ubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubKj	  )��}�(h�KCj  ]�h�j��  j  KubK j	  )��}�(h�KCj  ]�h�j��  j  K ubK!j	  )��}�(h�KCj  ]�h�j��  j  K!ubK"j	  )��}�(h�KCj  ]�h�j��  j  K"ubK#j	  )��}�(h�KCj  ]�h�j��  j  K#ubK$j	  )��}�(h�KCj  ]�h�j��  j  K$ubK%j	  )��}�(h�KCj  ]�h�j��  j  K%ubK&j	  )��}�(h�KCj  ]�h�j��  j  K&ubK'j	  )��}�(h�KCj  ]�h�j��  j  K'ubK(j	  )��}�(h�KCj  ]�h�j��  j  K(ubK)j	  )��}�(h�KCj  ]�h�j��  j  K)ubK*j	  )��}�(h�KCj  ]�h�j��  j  K*ubK+j	  )��}�(h�KCj  ]�h�j��  j  K+ubK,j	  )��}�(h�KCj  ]�h�j��  j  K,ubK-j	  )��}�(h�KCj  ]�h�j��  j  K-ubK.j	  )��}�(h�KCj  ]�h�j��  j  K.ubK/j	  )��}�(h�KCj  ]�h�j��  j  K/ubK0j	  )��}�(h�KCj  ]�h�j��  j  K0ubK1j	  )��}�(h�KCj  ]�h�j��  j  K1ubK2j	  )��}�(h�KCj  ]�h�j��  j  K2ubK3j	  )��}�(h�KCj  ]�h�j��  j  K3ubK4j	  )��}�(h�KCj  ]�h�j��  j  K4ubK5j	  )��}�(h�KCj  ]�h�j��  j  K5ubK6j	  )��}�(h�KCj  ]�h�j��  j  K6ubK7j	  )��}�(h�KCj  ]�h�j��  j  K7ubK8j	  )��}�(h�KCj  ]�h�j��  j  K8ubK9j	  )��}�(h�KCj  ]�h�j��  j  K9ubK:j	  )��}�(h�KCj  ]�h�j��  j  K:ubK;j	  )��}�(h�KCj  ]�h�j��  j  K;ubK<j	  )��}�(h�KCj  ]�h�j��  j  K<ubK=j	  )��}�(h�KCj  ]�h�j��  j  K=ubK>j	  )��}�(h�KCj  ]�h�j��  j  K>ubK?j	  )��}�(h�KCj  ]�h�j��  j  K?ubK@j	  )��}�(h�KCj  ]�h�j��  j  K@ubKAj	  )��}�(h�KCj  ]�h�j��  j  KAubKBj	  )��}�(h�KCj  ]�h�j��  j  KBubKCj	  )��}�(h�KCj  ]�h�j��  j  KCubuuj8  ]�j�8  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NKaK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKGKFKEKFKEKDKEKFKGKHKIKJKKKLKMKNKOKPKQKRKSKTKSKTKUKVKWKXKYKZK[K\K]K^K_K`KaKbNe]�(NK`K_K^K]NNKZKYKXKWKVKUKTKSKRKQKPKOKNNKLKKKJKIKHKGKFKEKFKEKDKEKDKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQKRKSKRKSKTKUKVKWKXNKZK[K\K]K^NK`KaNe]�(NK_K^K]K\K[NKYKXKWKVKUNNKRNKPKOKNKMKLKKNKIKHKGKFKEKDKEKDKCKDKCKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQKRKQKRKSKTKUKVKWKXKYKZK[K\K]K^K_K`Ne]�(NK^K]K\NKZKYKXKWNKUKTKSKRKQNKOKNKMKLKKKJKIKHKGKFKEKDKCKDKCKBKCKBKAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQKPKQKRKSKTKUKVKWKXKYKZK[K\K]K^K_Ne]�(NK]K\K[NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKCKBKAKBKAK@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKONKOKPNKTKSKTKUKVKWKXKYNK[K\K]K^Ne]�(NK\K[KZKYKXKWKVKUKTKSKRKQKPNKNKMKLKKKJKIKHKGKFKEKDKCKBKAKBKAK@KAK@K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNNKNKOKPNKRKSKTKUKVKWKXKYKZNK\K]Ne]�(NK[KZKYKXKWKVKUKTKSKRNKPKOKNKMKLKKNKINKGKFKEKDKCKBKAK@KAK@K?K@K?K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMNKMKNKOKPKQKRKSKTKUKVKWKXKYKZK[K\Ne]�(NKZKYNKWKVKUKTKSKRKQKPKONKMKLNKJKIKHKGKFKEKDKCKBKAK@K?K@K?K>K?K>K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKKKLKMNKOKPNKRKSKTKUKVKWKXKYKZK[Ne]�(NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKHNKDKCNNK@K?K>K?K>K=K>K=K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKJKKKLKMKNKONKQKRKSKTKUKVNKXKYKZNe]�(NKXKWKVKUKTKUKTNKPKOKNKMKLNKJKIKHKGKFNKDNKBKAK@K?K>K=NK=K<K=K<K;K<K=K>K?K@KAKBKCNKGKFKGKHKIKJKIKJKKKLKMKNKOKPKQKRNKTKUKVKWKXKYNe]�(NKWKVNKTKSKTNKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@NK>K=K<K=K<K;NNK:K;K<K=K>K?K@KAKBKCNKEKFKGKHKIKHKIKJKKKLKMKNKOKPNKRKSKTKUKVKWKXNe]�(NKVKUKTKSKRNKPKOKNKMKLKMNKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K<K;K:K9K:K9K:K;K<K=K>K?K@KAKBKCKDKEKFKGKHKGKHKIKJKKKLKMKNKOKPKQKRNKTKUKVKWNe]�(NKUKTKSKRKQKPKOKNNKLKKNKINKGKFKEKDKCKBKAK@NK>K=K<K;K:K;K:K9K8NK8K9K:K;K<K=K>K?K@KAKBKCKDNNKGKFKGKHKIKJKKKLKMKNKOKPKQKRKSKTKUKVNe]�(NKTKSKRKQKPKOKNKMKLKKKJNKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK9K8K7K8K7K8K9K:K;K<K=K>K?K@KANKCKDKEKFKEKFKGKHKIKJKKKLKMKNKOKPKQKRKSKTKUNe]�(NKSKRKQKPKOKNKMKLKKKJKIKHKGNKEKDKCKBKANK?K>K=K<K;K:K9K8NNK7K6NK6K7K8K9K:K;K<K=K>K?K@KAKBKCNKEKDKEKFKGKHKIKJKKNKOKNKOKPKQKRKSKTNe]�(NKRKQKPKOKNNKNNKJKIKHKGKFKEKDKCKBKAK@K?NK=K<K;NK9K8K7K6K7K6K5K6K5K6K7K8K9K:K;K<K=K>NK@KAKBKCKDKCKDKEKFKGKHKIKJNKNKMKNKOKPKQKRKSNe]�(NKQKPNKNKMKLKMKLKKKJNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K6K5K4K5K4K5K6K7K8K9K:K;K<K=K>K?K@KAKBNKBKCKDKEKFKGKHKIKJNKLKMKNKOKPKQKRNe]�(NKPKOKNKMKLKKKLKMKLKKNKEKDKCKBKCNK?K>K=K<K;NK9NK7NK5K4K5K4K3K4K3K4K5K6K7K8K9K:K;K<K=K>K?K@KAKBKAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQNe]�(NKOKNKMKLKKKJKKKLNNKENKCKBKANK?K>K=K<K;K:NK8K7K6K5NK3K4K3K2K3K2K3K4K5K6K7K8K9K:K;K<K=K>K?K@KAK@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPNe]�(NKNKMKLKKKJKINNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K3K2K1K2K1K2K3K4K5K6K7K8K9K:K;K<K=K>K?K@K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKONe]�(NKMKLKKNKIKHKGKFKENKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K2K1K0K1K0K1K2K3K4K5K6K7K8K9K:K;K<K=K>K?K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNNe]�(NKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0NK0K/NK/K0K1K2K3K4K5K6K7K8K9K:K;K<K=K>K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMNe]�(NKKKJKIKHNKFKENKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4K3NK1K0K/NK/K.K-K.K/K0K1K2K3K4K5K6K7K8K9K:K;K<K=K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLNe]�(NKJNKHKGKFNKDKCKBKCNK?K>K=K<K;K:K9K8NK6K5K4K3K2K1K0K/K.K/K.K-K,K-K.K/K0K1K2K3K4K5K6K7K8K9K:K;K<K;K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKNe]�(NKIKHKGKFKEKDKCKBKANK?K>K=K<K;K:K9K8K7NK5K4K3K2NK0K/NK-K.K-K,K+K,K-K.K/K0K1K2K3K4K5K6K7K8K9K:K;K:K;K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJNe]�(NKHKGKFKEKDKCKBKAK@K?NK=NNK:K9K8K7K6K5K4K3NK1K0K/K.K-K,K-K,K+K*NNNNNNNNNNNNNNNNK9K:K;K<K=K>K?K@NKDKCKDNKFKGKHKINe]�(NKGKFKEKDKCNKAK@K?K>K=K<K;K:K9K8NK6K5K4K3K2NK0K/K.K-K,K+K,K+K*K)NK+K,K-K.K/K0K1K2K3K4K5K6K7K8NK8K9K:K;K<K=K>K?K@NKBKCKDKEKFKGKHNe]�(NKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K1NK/K.K-K,K+K*K+K*K)K(NK*K+K,K-K.K/K0K1K2K3K4K5K6K7NK7K8K9K:K;K<K=K>K?K@KAKBKCKDKEKFKGNe]�(NKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7NK5K4K3K2K1K0K/K.K-K,K+K*K)K*K)K(K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6NK6K7K8K9K:K;K<K=K>K?K@KAKBKCKDKEKFNe]�(NKDKCKBKAK@NNNK<K;K:NK8NK6K5NK3K2K1K0K/K.K-K,K+K*K)K(K)K(K'K&NK*K+K,K-K.K/K0K1K2K3K4K5K6K7NK5K6K7K8K9K:K;K<NK>K?K@KAKBKCKDKENe]�(NKCKBKAK@K?K>NK<K;K:K9K8K7K6K5K4K3K2NK0K/K.K-K,K+K*K)K(K'K(K'K&K%NK+K,K-K.K/K0K1K2K3K4K5K6K7K8NK4K5K6K7K8K9K:K;K<K=K>K?K@KAKBKCKDNe]�(NKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-NK+K*K)K(K'K&K'K&K%K$NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NK3K4K5K6K7K8K9K:K;K<K=K>K?K@NKDKCNe]�(NKANK?K>NK<K;K:NK8K7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K&K%K$K#NNNNNNNNNNNNNNNNK2K3K4K5K6K7K8K9NK;K<K=K>NK@NKBNe]�(NK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K%NK#K"K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1NNK4K5K6K7K8NK:K;K<K=K>K?K@KANe]�(NK?NK=NK;K:K9K8K7NK5K4K3K2K1NK/K.K-K,K+K*K)K(K'NK%NK#NK#K"K!K K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4NK6K7NK9K:K;K<K=K>K?K@Ne]�(NK>K=K<K;K:NK8K7K6NK4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K#K"K!K KK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6NK8K9K:K;K<NK>K?Ne]�(NK=NNK:K9NK7K6K5K4K3NK1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K"K!K KKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2NK4K5K6K7K8K9K:K;K<K=K>Ne]�(NK<K;K:NK8K7K6K5K4K3K2K1K0K/K.K-K,NNK+NK'K&K%K$K#K"K!K K!K NKKKKK K!K"K#K$K%K&K'K(K)K*K+K,NK.K/K0K1K2K3K4NK6K7NNK:K;K<K=Ne]�(NK;K:K9K8K7K6K5K4K3K2K1K0K/K.NK,K+K*K)NNK&K%K$K#K"K!K KK KKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2NK4K5K6K7K8K9K:K;K<Ne]�(NK:K9K8K7K6K5K4K3K2NK0K/K.K-K,K+NK)K(K'K&K%NK#K"K!K KKNKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+NK-K.K/K0K1K2K3K4K5K6K7K8K9K:K;Ne]�(NK9K8K7K6K5NK3K2K1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!K NKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*NK,K-K.K/K0K1K2K3K4NK6K7K8K9K:Ne]�(NK8K7NK5K4K3K2K1K0K/K.K-K,NK*K)NK'K&K%K$K#K"K!K KKKKKKKNKKKKKNKNK!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7K8K9Ne]�(NK7K6K5K4K3K2NK0NK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKNKKK K!K"K#NK%K&NK(K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7K8Ne]�(NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K"NKKKNKKKKKKKKKKKKKNK K!K"K#K$K%K&K'K(NK*K+K,K-NK/K0K1K2K3K4K5K6K7Ne]�(NK5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$NK"K!K NKKKKKNKKKKKNNKNKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6Ne]�(NK4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#NK!K KNKKKKKKKNKKKKKKKNKKKKKK K!K"NK$K%K&K'K(NK*K+NK-K.K/K0K1K2K3K4K5Ne]�(NK3K2K1K0K/K.K-K,NK*K)K(K'NNNNK"K!K KKKKNKKKKKKKKKKKKKNKKKKKKK K!K"K#K$NK(K'K(K)K*K+K,K-K.K/K0K1K2K3K4Ne]�(NK2K1K0K/K.K-NK+NK)K(K'K&K%K$K#K"K!K KNKKKKNKKKNKKKKKKKKKKKKKKNKK K!NK#K$NK&K'K(NK*K+K,K-K.K/K0K1K2K3Ne]�(NK1K0K/K.NK,NK*K)K(K'K&K%K$K#K"K!K NKKKKKKKKKKNKKKKKKKKKKKKNKKKKK K!K"K#K$K%K&K'NK)K*K+K,K-K.K/K0K1K2Ne]�(NK0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKNKKKNKKKKKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1Ne]�(NK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKNKKKKKKKKKKKKKKKKNKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0Ne]�(NK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKNKKKKKKKKKKKKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/Ne]�(NK-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.Ne]�(NK,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKNKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-Ne]�(NK+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKNKKNKKKKKKKKKKKKKNKKNKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,Ne]�(NK*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKNKKKKKKKKKNKKKNKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+Ne]�(NK)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	K
KKKKKKKKKKKNKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*Ne]�(NK(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KNNNNNNNNKKKKKKKKKKKKKKKK K!K"K#K$K%K&K'K(K)Ne]�(NK'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKNK	K
KKKKNKKKKKKKKNKKNKKKKK K!K"K#K$K%K&K'K(Ne]�(NK&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKNKK	K
KKKNKKKKKKKKKKKNKKKKKK K!K"K#K$K%K&K'Ne]�(NK%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKKK	K
KKNKKKKKKKKKKKKNKKNKKK K!K"K#K$K%K&Ne]�(NK$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKNKK	K
KKKNKKKKKKKKNKKKKKKKKKKK K!K"K#K$K%Ne]�(NK#K"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKNK	K
KKKKNKKKKKKKKKKKKKNKKKKKKK K!K"K#K$Ne]�(NK"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKKNK
KKKKKNKKKKKKKKKKNKKKKKKKKKKK K!K"K#Ne]�(NK!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKKKK NNNNNNNK
KKKKKKKKKKKKKKKKKKKKKK K!K"Ne]�(NK"K!K KKKKKKKKKKKKKKKKKKKKKK
K	KKKKKKKKKKKKKKKK	K
KKKKKKKKKKKKKKKKKKKKKK K!Ne]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej�8  ]�j�8  aj�8  j�8  )��}�(j�8  ]�(�Player Ready: Kyle��
Game Start�ej�8  Kj�8  M�ubj�8  ]�h]aj�8  ]�(]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K KKK K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K KK K Ke]�(KK K K K K KK K K K K KKK KK K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K KK K K K KK K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K KK K K K Ke]�(KK K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K KK K K K K K K K K KK K Ke]�(KK K K K K K K K K K KK K K K K K KK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K Ke]�(KK K KK K K K K K K K K KK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K KK K KKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K Ke]�(KK K K K K K K KK K K K K KK K K K K KK KK K K K K K KK K K K K K K K K K K K K KK K K K K K K K K K K K K K K K KK K K K K K Ke]�(KK K KK K K KK K K K K K K K K K K K K K K K K KK K K K K K KKK K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K Ke]�(KK K K K K KK K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K Ke]�(KK K K K K K K K KK K KK KK K K K K K K K KK K K K K K K K K KK K K K K K K K K K K K K KKK K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K KK K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K KK K K K K KK K K K K K K K KKK K KK K K K K K K K K K K K K K KK K K K K K K K K KK K K K K K K K Ke]�(KK K K K K KK KK K K K K K K K K K K K KK K K KK K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K KK K K K K K K K Ke]�(KK K KK K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K KK K K K K K K Ke]�(KK K K K K K K K K K KK K K K K KK K K K K KK KK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K KKK KK K K KK K K K K K KK K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K KKK K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K KK K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K KK K KK K K K K K K K K K K KK K K K K KK K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK KK K K KK K K K KK K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K KK K K K K K K K K KK K K K KK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K KK KKK K K K K K K K KK K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K KK K K KK K K K Ke]�(KK K K K K KK K K K K K K K K K KK K K K K KK K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K KK K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K KK K K K KK K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K Ke]�(KK K K K K KKKK K K KK KK K KK K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K KK K K K K K K K Ke]�(KK K K K K K KK K K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K KK K Ke]�(KK KK K KK K K KK K K K K K K K K K K K K K KK K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K KK K K K KK KK Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K KKK K K K K KK K K K K K K K Ke]�(KK KK KK K K K K KK K K K K KK K K K K K K K K KK KK KK K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K Ke]�(KK K K K K KK K K KK K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K KK K Ke]�(KK KKK K KK K K K K KK K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K Ke]�(KK K K KK K K K K K K K K K K K K KKK KK K K K K K K K K K KK K K K K K K K K K K K K K K K K KK K K K K K K KK K KKK K K K Ke]�(KK K K K K K K K K K K K K K KK K K K KKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K Ke]�(KK K K K K K K K K KK K K K K K KK K K K K KK K K K K K KK K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K Ke]�(KK K K K K KK K K K K KK K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K KK K K K K Ke]�(KK K KK K K K K K K K K K KK K KK K K K K K K K K K K K K K K KK K K K K KK KK K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K KK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K KK K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K KK K K K K K KK K K KK K K K K K K K K K K K K KK K K K K K K K K KK K K K KK K K K K K K K K Ke]�(KK K K K K K K K K K K K K K KK K K KK K K KK K K K K KK K K K K KKK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K KK K K KK K K K K K K KK K K K K K K KK K K K K K K K KK K K K K KK K KK K K K K K K K K Ke]�(KK K K K K K K K KK K K K KKKKK K K K K K K KK K K K K K K K K K K K K KK K K K K K K K K K K KK K K K K K K K K K K K K K K Ke]�(KK K K K K K KK KK K K K K K K K K K K KK K K K KK K K KK K K K K K K K K K K K K K KK K K KK K KK K K KK K K K K K K K K K Ke]�(KK K K K KK KK K K K K K K K K K K KK K K K K K K K K K KK K K K K K K K K K K K KK K K K K K K K K K K K KK K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K KK K KK K K K K K K K K K K K K KK K KK K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K KK K K KK K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K KK K KK K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K K K K KK K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K K K K K K K KK K KK K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K KK K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K K K K K K KK K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KK K K K K K KK K K K K K K K K K KK K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K Ke]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKeej 9  ]�(j#9  j%9  j'9  j)9  j+9  j-9  ej.9  �Bricks
�j09  ]�(hj39  j59  j79  j99  j;9  j=9  j?9  jA9  jC9  hsjE9  jG9  jI9  jK9  jM9  jO9  eh{j��  jP9  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NK G�b      G�a�     G�a�     G�ap     G�a@     G�a     G�`�     G�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�L�     G�M@     G�N      G�M@     G�L�     Ne]�(NG�b      G�a�     G�a�     G�ap     NNG�`�     G�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     NG�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      NG�L�     G�K�     G�K      G�K�     G�L�     NG�L�     G�K�     Ne]�(NG�a�     G�a�     G�ap     G�a@     G�a     NG�`�     G�`�     G�`P     G�`      G�_�     NNG�^�     NG�^      G�]�     G�]@     G�\�     G�\�     G�\      NG�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�K      G�K�     G�L�     G�K�     G�K      Ne]�(NG�a�     G�ap     G�a@     NG�`�     G�`�     G�`�     G�`P     NG�_�     G�_�     G�_      G�^�     G�^`     NG�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�J@     G�K      G�K�     G�K      G�J@     Ne]�(NG�ap     G�a@     G�a     NG�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     NG�P      G�O�     NG�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     NG�J@     G�K      G�J@     G�I�     Ne]�(NG�a@     G�a     G�`�     G�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      NG�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     NG�O�     G�N�     G�N      NG�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�H�     G�I�     NG�I�     G�H�     Ne]�(NG�a     G�`�     G�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     NG�^      G�]�     G�]@     G�\�     G�\�     G�\      NG�[`     NG�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      NG�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�H      G�H�     G�H      G�H�     G�H      Ne]�(NG�`�     G�`�     NG�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     NG�\�     G�\�     NG�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     NG�K�     G�K      NG�I�     G�H�     G�H      G�G@     G�F�     G�G@     G�H      G�G@     G�H      G�G@     Ne]�(NG�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�[      NG�Y�     G�Y      NNG�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     NG�H�     G�H      G�G@     G�F�     G�E�     G�F�     NG�F�     G�G@     G�F�     Ne]�(NG�`�     G�`P     G�`      G�_�     G�_�     G�_�     G�_�     NG�^      G�]�     G�]@     G�\�     G�\�     NG�[�     G�[`     G�[      G�Z�     G�Z@     NG�Y�     NG�X�     G�X`     G�X      G�W�     G�W@     G�V�     NG�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     NG�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�H      NG�E      G�E�     G�E      G�E�     G�F�     G�E�     Ne]�(NG�`P     G�`      NG�_�     G�_      G�_�     NG�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      NG�W@     G�V�     G�V�     G�V      G�U�     G�U`     NNG�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     NG�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     NG�E      G�D@     G�E      G�D@     G�E      G�E�     G�E      Ne]�(NG�`      G�_�     G�_�     G�_      G�^�     NG�^      G�]�     G�]@     G�\�     G�\�     G�\�     NG�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     NG�C�     G�D@     G�E      G�D@     Ne]�(NG�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     NG�\�     G�\      NG�[`     NG�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      NG�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     NG�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      NNG�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�C�     G�B�     G�C�     G�D@     G�C�     Ne]�(NG�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     NG�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     NG�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     NG�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�B�     G�B      G�B�     G�C�     G�B�     Ne]�(NG�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     NG�Y�     G�Y�     G�Y      G�X�     G�X`     NG�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      NNG�S�     G�S�     NG�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     NG�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     NG�B�     G�B      G�A@     G�B      G�A@     G�B      G�B�     G�B      Ne]�(NG�^�     G�^`     G�^      G�]�     G�]@     NG�]@     NG�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     NG�V�     G�V�     G�V      NG�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      NG�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     NG�B      G�A@     G�@�     G�A@     G�@�     G�A@     G�B      G�A@     Ne]�(NG�^`     G�^      NG�]@     G�\�     G�\�     G�\�     G�\�     G�\      G�[�     NG�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     NG�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      NG�@�     G�?�     G�@�     G�?�     G�@�     G�A@     G�@�     Ne]�(NG�^      G�]�     G�]@     G�\�     G�\�     G�\      G�\�     G�\�     G�\�     G�\      NG�Y�     G�Y�     G�Y      G�X�     G�Y      NG�W�     G�W@     G�V�     G�V�     G�V      NG�U`     NG�T�     NG�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�?�     G�>      G�?�     G�@�     G�?�     Ne]�(NG�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�\      G�\�     NNG�Y�     NG�Y      G�X�     G�X`     NG�W�     G�W@     G�V�     G�V�     G�V      G�U�     NG�U      G�T�     G�T@     G�S�     NG�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�>      G�<�     G�>      G�?�     G�>      Ne]�(NG�]@     G�\�     G�\�     G�\      G�[�     G�[`     NNG�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     NG�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�<�     G�;      G�<�     G�>      G�<�     Ne]�(NG�\�     G�\�     G�\      NG�[`     G�[      G�Z�     G�Z@     G�Y�     NG�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�;      G�9�     G�;      G�<�     G�;      Ne]�(NG�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      NG�Q@     G�P�     NG�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�9�     G�8      G�9�     G�;      G�9�     Ne]�(NG�\�     G�\�     G�\      G�[�     NG�[      G�Z�     NG�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      NG�T�     G�T@     G�S�     G�S�     G�S      NG�R`     G�R      G�Q�     NG�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�8      G�6�     G�8      G�9�     G�8      Ne]�(NG�\�     NG�[�     G�[`     G�[      NG�Z@     G�Y�     G�Y�     G�Y�     NG�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     NG�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�6�     G�5      G�6�     G�8      G�6�     Ne]�(NG�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      NG�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     NG�T�     G�T@     G�S�     G�S�     NG�R�     G�R`     NG�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�5      G�3�     G�5      G�6�     G�5      Ne]�(NG�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     NG�W�     NNG�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     NG�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     NNNNNNNNNNNNNNNNG�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      NG�5      G�3�     G�2      NG�2      G�3�     G�5      G�3�     Ne]�(NG�[`     G�[      G�Z�     G�Z@     G�Y�     NG�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     NG�U      G�T�     G�T@     G�S�     G�S�     NG�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     NG�P      G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      G�S�     G�S�     G�T@     G�T�     G�U      NG�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      NG�2      G�0�     G�.      G�0�     G�2      G�3�     G�2      Ne]�(NG�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      NG�T@     G�S�     G�S�     G�S      NG�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      NG�O�     G�P      G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      G�S�     G�S�     G�T@     G�T�     NG�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�.      G�0�     G�2      G�0�     Ne]�(NG�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     NG�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�N      G�N�     G�O�     G�P      G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      G�S�     G�S�     G�T@     NG�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�(      G�+      G�.      G�0�     G�.      Ne]�(NG�Z@     G�Y�     G�Y�     G�Y      G�X�     NNNG�W@     G�V�     G�V�     NG�U�     NG�U      G�T�     NG�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     NG�O�     G�P      G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      G�S�     G�S�     G�T@     G�T�     NG�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      NG�.      G�+      G�(      G�%      G�(      G�+      G�.      G�+      Ne]�(NG�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      NG�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     NG�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     NG�P      G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      G�S�     G�S�     G�T@     G�T�     G�U      NG�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�(      G�%      G�"      G�%      G�(      G�+      G�(      Ne]�(NG�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     NG�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      NG�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      G�S�     G�S�     G�T@     G�T�     G�U      G�U`     NG�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�(      G�%      G�"      G�      G�"      NG�(      G�%      Ne]�(NG�Y      NG�X`     G�X      NG�W@     G�V�     G�V�     NG�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     NG�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     NNNNNNNNNNNNNNNNG�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     NG�%      G�"      G�      G�      NG�      NG�"      Ne]�(NG�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�M@     NG�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     NNG�5      G�3�     G�2      G�0�     G�.      NG�"      G�      G�      G�      G�      G�      G�      G�      Ne]�(NG�Y      NG�X`     NG�W�     G�W@     G�V�     G�V�     G�V      NG�U`     G�U      G�T�     G�T@     G�S�     NG�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     NG�M@     NG�K�     NG�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      NG�.      G�+      NG�      G�      G�      G�      G��      G�      G�      G�      Ne]�(NG�Y�     G�Y      G�X�     G�X`     G�X      NG�W@     G�V�     G�V�     NG�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     NG�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�(      NG�      G�      G�      G��      G�       NG�      G�      Ne]�(NG�Y�     NNG�X      G�W�     �      NG�V�     G�V�     G�V      G�U�     G�U`     NG�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     NG�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      NG�(      G�%      G�"      G�      G�      G�      G�      G��      G�      G�      G�      Ne]�(NG�Y�     G�Y      G�X�     NG�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     NNG�Q�     NG�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      NG�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      NG�5      G�3�     G�2      G�0�     G�.      G�+      G�(      NG�"      G�      NNG�      G�      G�      G�      Ne]�(NG�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     NG�S�     G�S      G�R�     G�R`     NNG�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      NG�(      G�%      G�"      G�      G�      G�      G�      G�      G�"      Ne]�(NG�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     NG�U�     G�U`     G�U      G�T�     G�T@     G�S�     NG�R`     G�R      G�Q�     G�Q@     G�P�     NG�P      G�O�     G�N�     G�N      G�M@     G�L�     NG�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     NG�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�(      G�%      G�"      G�      G�      G�      G�"      G�%      Ne]�(NG�Y�     G�Y�     G�Y      G�X�     G�X`     NG�W�     G�W@     G�V�     G�V�     G�V      NG�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     NG�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      NG�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�(      NG�"      G�      G�"      G�%      G�(      Ne]�(NG�Z@     G�Y�     NG�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      NG�T@     G�S�     NG�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     NG�J@     G�I�     G�H�     G�H      G�G@     NG�E�     NG�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�(      G�%      G�"      G�%      G�(      G�+      Ne]�(NG�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      NG�W@     NG�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      NG�F�     G�E�     G�E      G�D@     G�C�     G�B�     NG�A@     G�@�     NG�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�(      G�%      G�(      G�+      G�.      Ne]�(NG�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     NG�S�     G�S�     G�S      G�R�     G�R`     G�R      NG�Q@     G�P�     G�P�     NG�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     NG�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      NG�;      G�9�     G�8      G�6�     NG�3�     G�2      G�0�     G�.      G�+      G�(      G�+      G�.      G�0�     Ne]�(NG�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     NG�U      G�T�     G�T@     NG�S�     G�S      G�R�     NG�R      G�Q�     G�Q@     G�P�     G�Q@     NG�O�     G�N�     G�N      G�M@     G�L�     NNG�J@     NG�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�.      G�0�     G�2      Ne]�(NG�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     NG�S�     G�S�     G�S      NG�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      NG�N�     G�N      G�M@     G�L�     G�K�     G�K      G�K�     NG�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     NG�B      G�A@     G�@�     G�?�     G�>      NG�;      G�9�     NG�6�     G�5      G�3�     G�2      G�0�     G�.      G�0�     G�2      G�3�     Ne]�(NG�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     NG�X      G�W�     G�W@     G�V�     NNNNG�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     NG�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�L�     NG�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      NG�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�2      G�3�     G�5      Ne]�(NG�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     NG�Y      NG�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     NG�S�     G�S�     G�S      G�S�     NG�R      G�Q�     G�Q@     NG�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     NG�E�     G�E      G�D@     NG�B�     G�C�     NG�@�     G�?�     G�>      NG�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�3�     G�5      G�6�     Ne]�(NG�\      G�[�     G�[`     G�[      NG�Z@     NG�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     NG�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     NG�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     NG�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     NG�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�5      G�6�     G�8      Ne]�(NG�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     NG�R      G�Q�     G�Q@     NG�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�6�     G�8      G�9�     Ne]�(NG�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      NG�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     NG�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�8      G�9�     G�;      Ne]�(NG�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     NG�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�9�     G�;      G�<�     Ne]�(NG�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�;      G�<�     G�>      Ne]�(NG�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     NG�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�<�     G�>      G�?�     Ne]�(NG�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      NG�T@     G�S�     NG�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     NG�K�     G�K      NG�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�>      G�?�     G�@�     Ne]�(NG�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      NG�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     NG�M@     G�L�     G�K�     NG�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�>      G�?�     G�@�     G�A@     Ne]�(NG�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     NG�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�?�     G�@�     G�A@     G�B      Ne]�(NG�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     NNNNNNNNG�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�@�     G�A@     G�B      G�B�     Ne]�(NG�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     NG�V      G�V�     G�V�     G�W@     G�W�     G�X      NG�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     NG�J@     G�I�     NG�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�A@     G�B      G�B�     G�C�     Ne]�(NG�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     NG�U�     G�V      G�V�     G�V�     G�W@     G�W�     NG�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     NG�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�B      G�B�     G�C�     G�D@     Ne]�(NG�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�U      G�U`     G�U�     G�V      G�V�     G�V�     G�W@     NG�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�K�     NG�H�     G�H      NG�F�     G�E�     G�E      G�D@     G�C�     G�B�     G�C�     G�D@     G�E      Ne]�(NG�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      NG�U�     G�V      G�V�     G�V�     G�W@     G�W�     NG�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      NG�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     G�D@     G�E      G�E�     Ne]�(NG�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     NG�V      G�V�     G�V�     G�W@     G�W�     G�X      NG�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      NG�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�E      G�E�     G�F�     Ne]�(NG�`�     G�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     NG�V�     G�V�     G�W@     G�W�     G�X      G�X`     NG�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      NG�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�E�     G�F�     G�G@     Ne]�(NG�a     G�`�     G�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�V�     NNNNNNNG�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�F�     G�G@     G�H      Ne]�(NG�a@     G�a     G�`�     G�`�     G�`�     G�`P     G�`      G�_�     G�_�     G�_      G�^�     G�^`     G�^      G�]�     G�]@     G�\�     G�\�     G�\      G�[�     G�[`     G�[      G�Z�     G�Z@     G�Y�     G�Y�     G�Y      G�X�     G�X`     G�X      G�W�     G�W@     G�V�     G�V�     G�V      G�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�O�     G�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�G@     G�H      G�H�     Ne]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej�9  j��  j��  M�j��  �ground, covered in leaves
�j��  ]�(]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  h"j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  haj��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j́  j��  j��  j��  j��  j��  j��  j��  j��  j΁  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  h"j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jс  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jՁ  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  haj��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jс  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j΁  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  haj��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j́  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jс  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  h"j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  haj��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  j��  jс  j��  j��  j��  j��  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  jɁ  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  e]�(j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  j��  eej��  j��  j��  ]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKK KKKKKK K K KK e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K KK e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K KK e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K KK Ke]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK KKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K KKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKK K K K KKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKK K K K K KKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K eej?�  ]�(KKejA�  ]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKK KKK K K KKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K KK e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K KKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK KKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK KKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK KKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKK KKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K KKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K K KKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKK K KKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKK K K K KKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKe]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K eej�9  hj��  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NKaK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K&K%K$K#K"Ne]�(NK`K_K^K]NNKZKYKXKWKVKUKTKSKRKQKPKOKNNKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K%K$NK"K!Ne]�(NK_K^K]K\K[NKYKXKWKVKUNNKRNKPKOKNKMKLKKNKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K$K#K"K!K Ne]�(NK^K]K\NKZKYKXKWNKUKTKSKRKQNKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K#K"K!K KNe]�(NK]K\K[NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-NK+K*NK(K'K&K%K$K#K"K!NK!K KKNe]�(NK\K[KZKYKXKWKVKUKTKSKRKQKPNKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,NK*K)K(NK&K%K$K#K"K!K K!K NKKNe]�(NK[KZKYKXKWKVKUKTKSKRNKPKOKNKMKLKKNKINKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K!K KK KKKKNe]�(NKZKYNKWKVKUKTKSKRKQKPKONKMKLNKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$NK"K!K KKKKKKKNe]�(NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKHNKDKCNNK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#NK!K KKKKNKKKNe]�(NKXKWKVKUKTKUKTNKPKOKNKMKLNKJKIKHKGKFNKDNKBKAK@K?K>K=NK;K:K9K8K7K6K5K4K3K2K1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!K KK NKKKKKKNe]�(NKWKVNKTKSKTNKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@NK>K=K<K;K:K9NNK6K5K4K3K2K1K0K/K.K-NK+K*K)K(K'K&K%K$K#K"K!K KKNKKKKKKKNe]�(NKVKUKTKSKRNKPKOKNKMKLKMNKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKNKKKKNe]�(NKUKTKSKRKQKPKOKNNKLKKNKINKGKFKEKDKCKBKAK@NK>K=K<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+K*K)K(NNK%K$K#K"K!K KKKKKKKKKKKKNe]�(NKTKSKRKQKPKOKNKMKLKKKJNKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4K3K2K1K0K/K.K-K,K+K*K)NK'K&K%K$K#K"K!K KKKKKKKKKKKKKNe]�(NKSKRKQKPKOKNKMKLKKKJKIKHKGNKEKDKCKBKANK?K>K=K<K;K:K9K8NNK5K4NK2K1K0K/K.K-K,K+K*K)K(K'K&K%NK#K"K!K KKKKKNKKKKKKKKNe]�(NKRKQKPKOKNNKNNKJKIKHKGKFKEKDKCKBKAK@K?NK=K<K;NK9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K KKKKKKNKKKKKKKKNe]�(NKQKPNKNKMKLKMKLKKKJNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"NK KKKKKKKKNKKKKKKKNe]�(NKPKOKNKMKLKKKLKMKLKKNKEKDKCKBKCNK?K>K=K<K;NK9NK7NK5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKNe]�(NKOKNKMKLKKKJKKKLNNKENKCKBKANK?K>K=K<K;K:NK8K7K6K5NK3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKNe]�(NKNKMKLKKKJKINNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKNe]�(NKMKLKKNKIKHKGKFKENKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKNe]�(NKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0NK.K-NK+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKNe]�(NKMKLKKKJNKHKGNKEKDKCKBKAK@K?K>K=K<K;NK7K6K5K4K3NK1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKNe]�(NKNNKLKKKJNKHKGKFKENKCKBKAK@K?K>K=K<NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKNe]�(NKMKLKKKJKIKHKGKFKENKCKBKAK@K?K>K=K<K;NK7K6K5K4NK2K1NK-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKK
Ne]�(NKLKKKJKIKHKGKFKEKDKCNKANNK>K=K<K;K:K9K8K7NK3K2K1K0K/K.K-K,K+K*NNNNNNNNNNNNNNNNKKKKKKKKNKKKNKKK
K	Ne]�(NKKKJKIKHKGNKEKDKCKBKAK@K?K>K=K<NK:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+NK-K.K/K0K1K2K3K4K5K6K7K8K9K:NKKKKKKKKKNKKK
KK
K	KNe]�(NKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK8K7K6K5NK3K2K1K0K/K.K-K,K+K*NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NKKKKKKKKKKKK
K	K
K	KKNe]�(NKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=NK9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7K8NKKKKKKKKKKK
K	KK	KKKNe]�(NKJKIKHKGKFNNNKBKAK@NK>NK<K;NK7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NKKKKKKKKNK
K	KKKKKKNe]�(NKIKHKGKFKEKDNKBKAK@K?K>K=K<K;K:K9K8NK4K3K2K1K0K/K.K-K,K+K*K)K(K'NK-K.K/K0K1K2K3K4K5K6K7K8K9K:NKKKKKKKKK
K	KKKKKKKNe]�(NKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3NK/K.K-K,K+K*K)K(K'K&NK.K/K0K1K2K3K4K5K6K7K8K9K:K;NKKKKKKKK
K	KKKKKNKKNe]�(NKGNKEKDNKBKAK@NK>K=K<K;K:K9K8K7K6K5K4K3K2K1NK-K,K+K*K)K(K'K&K%NNNNNNNNNNNNNNNNKKKKKKKKNKKKKNKNKNe]�(NKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)NK%K$K#K"K!K KKKKKKKKKKKKKNNKKKKKNKKKKKKK KNe]�(NKGNKENKCKBKAK@K?NK=K<K;K:K9NK5K4K3K2K1K0K/K.K-NK+NK)NK'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKNKKNKKKKKKKKNe]�(NKHKGKFKEKDNKBKAK@NK<K;K:K9K8K7K6K5K4K3NK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKNKKKKKNKKNe]�(NKINNKDKCNKAK@K?K>K=NK9K8K7K6K5K4K3K2K1K0NK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKNKKK
K	KKKKKKKNe]�(NKHKGKFNKBKAK@K?K>K=K<K;K:K9K8K7K6NNK3NK1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K KKKKKKKKKKNKKKKKKKNK
K	NNKKKKNe]�(NKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK8K7K6K5NNK0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKNKKK
K	KKKKKNe]�(NKHKGKFKEKDKCKBKAK@NK>K=K<K;K:K9NK5K4K3K2K1NK/K.K-K,K+K*NK(K'K&K%K$K#K"K!K KKKKKKKKKKKNKKKKKKKKKK
K	KKKKNe]�(NKIKHKGKFKENKCKBKAK@K?NK;K:K9K8K7K6K5K4K3K2K1K0K/K.NK,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKNKKKKKKKKKNK
K	KKKNe]�(NKJKINKEKDKCKBKAK@K?K>K=K<NK:K9NK7K6K5K4K3K2K1K0K/K.K-K,K+K*K)NK'K&K%K$K#NK!NKKKKKKKKKKKKKKKKKKKKKK
K	KK	Ne]�(NKIKHKGKFKEKDNKBNK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$NK"K!K KKKNKKNKKKKKKKKKKKKKKK
K	K
Ne]�(NKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;NK9K8K7K6K5K4NK2K1K0NK.K-K,K+K*K)K(K'K&K%K$K#K"NK KKKKKKKKNKKKKNKKKKKKKK
KNe]�(NKKKJKIKHKGKFKEKDKCKBKAK@K?K>NK<K;K:NK8K7K6NK4K3K2K1K2NK.K-K,K+K*NNK'NK%K$K#K"K!K KKKKKKKKKKKKKKKKKK�      KKKKNe]�(NKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;NK9K8K7NK5K4K3K2K1K0K/NK-K,K+K*K)K(K)NK%K$K#K"K!K KKNKKKKKNKKNKKKKKKKKKNe]�(NKMKLKKKJKIKHKGKFNKDKCKBKANNNNK<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+K*K)K*NK&K%K$K#K"K!K KKKKNKKKKKKKKKKKKKKKNe]�(NKNKMKLKKKJKINKGNKEKDKCKBKAK@K?K>K=K<K;NK9K8K7K8NK4K3K2NK0K/K.K-K,K+K*K)K(K'K&K%K$K#NK!K KNKKNKKKNKKKKKKKKKKNe]�(NKOKNKMKLNKJNKHKGKFKEKDKCKBKAK@K?K>NK<K;K:K9K8K7K6K5K4K3NK1K0K/K.K-K,K+K*K)K(K'K&NK$K#K"K!K KKKKKKKNKKKKKKKKKKNe]�(NKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2NK0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKNe]�(NKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7NK5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&NK$K#K"K!K KKKKKKKKKKKKKKKKNe]�(NKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKNe]�(NKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKNe]�(NKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*NK(K'K&K%K$K#K"K!K KKKKKKKKKKKKKNe]�(NKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NK:K9NK7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(NK&K%K$K#K"K!K KKKKKKKKKKKKNe]�(NKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7NK5K4K3K2K1K0K/K.K-NK+K*K)NK'K&K%K$K#K"K!K KKKKKKKKKKKNe]�(NKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K!K KKKKKKKKKKNe]�(NKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8NNNNNNNNK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKNe]�(NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK?K@KAKBKCKDNK0K/K.K-K,K+K*K)NK'K&NK$K#K"K!K KKKKKKKKNe]�(NKZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK>K?K@KAKBKCNK1K0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K KKKKKKKNe]�(NK[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K<K=K>K?K@KAKBNK2K1K0K/K.K-K,K+K*K)K(K)NK%K$NK"K!K KKKKKKNe]�(NK\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NK>K?K@KAKBKCNK3K2K1K0K/K.K-K,NK*K)K(K'K&K%K$K#K"K!K KKKKKNe]�(NK]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=NK?K@KAKBKCKDNK4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K KKKKNe]�(NK^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>NK@KAKBKCKDKENK5K4K3K2K1K0K/K.K-K,NK*K)K(K'K&K%K$K#K"K!K KKKNe]�(NK_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K@NNNNNNNK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KK Ne]�(NK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K K!Ne]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej͂  ]�(K"KAejς  ]�(h]j҂  jԂ  jւ  j؂  hj39  j59  j79  j99  j;9  j=9  j?9  jA9  jC9  hsjE9  jG9  jI9  jK9  jM9  jO9  ej  }�(K h})��}�(h�Kh�K h!h"h�j��  j  K'h&�Item�h|j=9  )��}�(h{j�  hKhKhKhj��  hj��  h�h�hKh �h!h"h#Kh$�h%Kh&�Bow�h(�ububKh})��}�(h�Kh�Kh!j��  h�j��  j  K#h&�Enemy�h|j'9  )��}�(hK
hK hj=9  )��}�(hKhKhKhj��  hj��  h�h�hKh �h!h"h#Kh$�h%Kh&j�  h(�ubhKh)�h*�j�  �h+Kh,�h!j��  h7K	hKh8K hK hphs)��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j��  hj��  ubj�  G?�      hfKhNNj�  Nhn]�hPKdhRKh&�Goblin Archer�hTK hY]�hMK hg]�h]�(K�KKej�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&�Leather Shirt�hjƄ  ubj��  ]�(j�  h})��}�(h�Kh�Kh!j��  h�j��  j  K'h&j�  h|j)9  )��}�(hKhK hj99  )��}�(hKhKhKhj��  h�1H�h�h�hKh �h!h"h#Kh$�h%Kh&�	Longsword�h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjK9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&�	Iron Helm�hj��  ubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&�Goblin Knight�hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j�  hjƄ  ubj��  ]�(j�  j�  ej�  j79  )��}�(hKhKhj��  hj%�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&�Wooden Shield�hK ubj�  �h%Kububej�  Nj�  �h%KububKj�  Kh})��}�(h�Kh�Kh!j��  h�j��  j  K8h&j�  h|j+9  )��}�(hK	hK hj99  )��}�(hKhKhKhj��  hj%�  h�h�hKh �h!h"h#Kh$�h%Kh&j&�  h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hj��  h&�Leather Helm�hj��  ubj�  G?��Q�hfKhNNj�  Nhn]�hPKdhRKh&�Goblin Grunt�hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j4�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j�  hjƄ  ubj��  ]�(j4�  h})��}�(h�Kh�Kh!j��  h�j��  j  K6h&j�  h|j%9  )��}�(hKhK hj;9  )��}�(hKhKhKhj��  hj��  h�h�hKh �h!h"h#Kh$�h%Kh&�
Greatsword�h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hj��  h&j<�  hj��  ubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&�Goblin Berserker�hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{jD�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j�  hjƄ  ubj��  ]�(j4�  jD�  ej�  Nj�  �h%Kububej�  Nj�  �h%KububKh})��}�(h�Kh�Kh!hah�j��  j  K5h&�Health�h|h])��}�(h`Kh�h(�h!hah{jT�  hj��  h&j��  hj��  ububKjD�  Kh})��}�(h�Kh�Kh!j��  h�j��  j  K(h&j�  h|j'9  )��}�(hK
hK hj=9  )��}�(hKhKhKhj��  hj��  h�h�hKh �h!h"h#Kh$�h%Kh&j�  h(�ubhKh)�h*�j�  �h+Kh,�h!j��  h7KhKh8K hK hphs)��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j��  hj��  ubj�  G?�      hfKhNNj�  Nhn]�hPKdhRKh&j�  hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{jY�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j�  hjƄ  ubj��  ]�(jY�  h})��}�(h�Kh�Kh!j��  h�j��  j  K+h&j�  h|j#9  )��}�(hK	hK hj?9  )��}�(hKhKhKhj��  hj��  h�h�hKh �h!h"h#Kh$�h%Kh&�Spear�h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hj��  h&j<�  hj��  ubj�  G?�������hfKhNNj�  Nhn]�hPKdhRKh&�Goblin Lancer�hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{jg�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j�  hjƄ  ubj��  ]�(jY�  jg�  h})��}�(h�Kh�K
h!j��  h�j��  j  K#h&j�  h|j%9  )��}�(hKhK hj;9  )��}�(hKhKhKhj��  hj��  h�h�hKh �h!h"h#Kh$�h%Kh&jJ�  h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hj��  h&j<�  hj��  ubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&jN�  hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{jw�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j�  hjƄ  ubj��  ]�(jY�  jw�  ej�  Nj�  �h%Kububh})��}�(h�Kh�Kh!jс  h�j��  j  K.h&j�  h|j�8  )��}�(hKhK hjj�  )��}�(hKhKhKhj��  hj%�  h�h�hKh �h!h"h#Kh$�h%Kh&�Mace�h(�ubhKh)�h*�j�  �h+K h,�h!jс  h7K	hKh8K hK hpjK9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j)�  hj��  ubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&�Goblin Stonewall�hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j��  j��  jI9  )��}�(h�h(�hKh!h"h#K7h8K2h$�hj��  h&�Iron Breastplate�hjƄ  ubj��  ]�(jg�  j��  ej�  j39  )��}�(hKhKhj��  hj%�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&�Iron Shield�hK ubj�  �h%Kububej�  j59  )��}�(hKhKhj��  hjɄ  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&�Buckler�hK ubj�  �h%Kububjw�  j��  ej�  Nj�  �h%KububKjg�  Kh})��}�(h�Kh�Kh!j΁  h�j��  j  K+h&�Chest�h|j��  )��}�(h{j��  hY]�(jM9  )��}�(h�h(�hKh!h"h#K#h8K#h$�hj��  h&�Chain Shirt�hjƄ  ubjA9  )��}�(hKhKhKhj��  hj%�  h�h�hKh �h!h"h#Kh$�h%Kh&�Dagger�h(�ubj79  )��}�(hKhKhj��  hj%�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&j3�  hK ubj��  )��}�(h�j��  Kh(�h!j��  h]�(K�K�Keh&�
Gold Coins�hj��  ubeh!j΁  h]�(KQKOKeh&j��  ububK	h})��}�(h�Kh�K	h!h"h�j��  j  K(h&j	�  h|j79  )��}�(h{j��  hKhKhj��  hj%�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&j3�  hK ububK
jw�  Kj��  Kh})��}�(h�K"h�Kh!jՁ  h�j��  j  KAh&�	Stairs Up�h|j��  )��}�(h{j��  h�K"h�J����h�j��  j  KAj��  Kh&�Stairs�h|NububKj��  Kh})��}�(h�K5h�Kh!hah�j��  j  K=h&jV�  h|h])��}�(h`Kh�h(�h!hah{j��  hj��  h&j��  hj��  ububKh})��}�(h�K7h�Kh!jс  h�j��  j  K=h&j�  h|j�8  )��}�(hKhK hjj�  )��}�(hKhKhKhj��  hj%�  h�h�hKh �h!h"h#Kh$�h%Kh&j��  h(�ubhKh)�h*�j�  �h+K h,�h!jс  h7KhKh8K hK hpjK9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j)�  hj��  ubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&j��  hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j��  j��  jI9  )��}�(h�h(�hKh!h"h#K7h8K2h$�hj��  h&j��  hjƄ  ubj��  ]�(j��  h})��}�(h�K7h�Kh!j��  h�j��  j  K@h&j�  h|j%9  )��}�(hKhK hj;9  )��}�(hKhKhKhj��  hj��  h�h�hKh �h!h"h#Kh$�h%Kh&jJ�  h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hj��  h&j<�  hj��  ubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&jN�  hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j˿  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j�  hjƄ  ubj��  ]�(j��  j˿  ej�  Nj�  �h%Kububej�  j39  )��}�(hKhKhj��  hj%�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&j��  hK ubj�  �h%KububKj˿  Kh})��}�(h�K;h�Kh!j΁  h�j��  j  Kh&j��  h|j��  )��}�(h{jۿ  hY]�(j39  )��}�(hKhKhj��  hj%�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&j��  hK ubj39  )��}�(hKhKhj��  hj%�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&j��  hK ubhs)��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j��  hj��  ubj��  )��}�(h�j��  Kh(�h!j��  hj��  h&j��  hj��  ubeh!j΁  hj��  h&j��  ububKh})��}�(h�K<h�Kh!j��  h�j��  j  Kh&j�  h|j%9  )��}�(hKhK hj;9  )��}�(hKhKhKhj��  hj��  h�h�hKh �h!h"h#Kh$�h%Kh&jJ�  h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hj��  h&j<�  hj��  ubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&jN�  hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j�  hjƄ  ubj��  ]�(j�  h})��}�(h�K>h�Kh!jс  h�j��  j  Kh&j�  h|j�8  )��}�(hKhK hjj�  )��}�(hKhKhKhj��  hj%�  h�h�hKh �h!h"h#Kh$�h%Kh&j��  h(�ubhKh)�h*�j�  �h+K h,�h!jс  h7KhKh8K hK hpjK9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j)�  hj��  ubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&j��  hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j��  j��  jI9  )��}�(h�h(�hKh!h"h#K7h8K2h$�hj��  h&j��  hjƄ  ubj��  ]�(j�  j��  ej�  j39  )��}�(hKhKhj��  hj%�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&j��  hK ubj�  �h%Kububej�  Nj�  �h%KububKh})��}�(h�K=h�Kh!j��  h�j��  j  Kh&j�  h|j+9  )��}�(hK	hK hj99  )��}�(hKhKhKhj��  hj%�  h�h�hKh �h!h"h#Kh$�h%Kh&j&�  h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hj��  h&j<�  hj��  ubj�  G?��Q�hfKhNNj�  Nhn]�hPKdhRKh&j>�  hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j�  hjƄ  ubj��  ]�(j�  h})��}�(h�K=h�Kh!j��  h�j��  j  Kh&j�  h|j'9  )��}�(hK
hK hj=9  )��}�(hKhKhKhj��  hj��  h�h�hKh �h!h"h#Kh$�h%Kh&j�  h(�ubhKh)�h*�j�  �h+Kh,�h!j��  h7KhKh8K hK hphs)��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j��  hj��  ubj�  G?�      hfKhNNj�  Nhn]�hPKdhRKh&j�  hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j�  hjƄ  ubj��  ]�(j�  j�  j�  h})��}�(h�K>h�Kh!j��  h�j��  j  Kh&j�  h|j'9  )��}�(hK
hK hj=9  )��}�(hKhKhKhj��  hj��  h�h�hKh �h!h"h#Kh$�h%Kh&j�  h(�ubhKh)�h*�j�  �h+Kh,�h!j��  h7KhKh8K hK hphs)��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j��  hj��  ubj�  G?�      hfKhNNj�  Nhn]�hPKdhRKh&j�  hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j"�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j�  hjƄ  ubj��  ]�(j�  j�  j"�  ej�  Nj�  �h%Kububej�  Nj�  �h%Kububj"�  ej�  Nj�  �h%KububKj�  Kh})��}�(h�K=h�Kh!hah�j��  j  Kh&jV�  h|h])��}�(h`Kh�h(�h!hah{j0�  hj��  h&j��  hj��  ububKj"�  Kj��  Kh})��}�(h�K?h�Kh!h"h�j��  j  Kh&j	�  h|j59  )��}�(h{j4�  hKhKhj��  hjɄ  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&j��  hK ububKh})��}�(h�K?h�Kh!hah�j��  j  K'h&jV�  h|h])��}�(h`Kh�h(�h!hah{j8�  hj��  h&j��  hj��  ububKh})��}�(h�K@h�Kh!jс  h�j��  j  K$h&j�  h|j�8  )��}�(hKhK hjj�  )��}�(hKhKhKhj��  hj%�  h�h�hKh �h!h"h#Kh$�h%Kh&j��  h(�ubhKh)�h*�j�  �h+K h,�h!jс  h7K	hKh8K hK hpjK9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j)�  hj��  ubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&j��  hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{j<�  j��  jI9  )��}�(h�h(�hKh!h"h#K7h8K2h$�hj��  h&j��  hjƄ  ubj��  ]�(j<�  h})��}�(h�K@h�Kh!j��  h�j��  j  K%h&j�  h|j%9  )��}�(hKhK hj;9  )��}�(hKhKhKhj��  hj��  h�h�hKh �h!h"h#Kh$�h%Kh&jJ�  h(�ubhKh)�h*�j�  �h+K h,�h!j��  h7KhKh8K hK hpjG9  )��}�(h�h(�hKh!h"h#Kh8K
h$�hj��  h&j<�  hj��  ubj�  G        hfKhNNj�  Nhn]�hPKdhRKh&jN�  hTK hY]�hMK hg]�hj�  j�  NhjK j�  K(j�  K j�  NhO�hmNhxKhy�j��  Kh{jJ�  j��  jE9  )��}�(h�h(�hKh!h"h#Kh8Kh$�hj��  h&j�  hjƄ  ubj��  ]�(j<�  jJ�  ej�  Nj�  �h%Kububej�  j39  )��}�(hKhKhj��  hj%�  h�h�h(�h �h!h"h#Kh8Kh$�h%K h&j��  hK ubj�  �h%KububKjJ�  Kh})��}�(h�KAh�Kh!j��  h�j��  j  K"h&�Stairs Down�h|jL�  )��}�(h{jZ�  h|Nh�J����h�j��  h�KAj��  Kh&j��  j  K"ububujO�  ]�(h]j҂  jԂ  jւ  j؂  eh&�
1B: Forest�jR�  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NK`K_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K%K$K#K"K!Ne]�(NK_K^K]K\NNKYKXKWKVKUKTKSKRKQKPKOKNKMNKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$K#K$K#NK!K Ne]�(NK^K]K\K[KZNKXKWKVKUKTNNKQNKOKNKMKLKKKJNKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K#K"K!K KNe]�(NK]K\K[NKYKXKWKVNKTKSKRKQKPNKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K"K!K KKNe]�(NK\K[KZNKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,NK*K)NK'K&K%K$K#K"K!K NK KKKNe]�(NK[KZKYKXKWKVKUKTKSKRKQKPKONKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+NK)K(K'NK%K$K#K"K!K KK KNKKNe]�(NKZKYKXKWKVKUKTKSKRKQNKOKNKMKLKKKJNKHNKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*NK(K'K&K%K$K#K"K!K KKKKKKKNe]�(NKYKXNKVKUKTKSKRKQKPKOKNNKLKKNKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&NK$K#NK!K KKKKKKKKNe]�(NKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKGNKCKBNNK?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"NK KKKKKNKKKNe]�(NKWKVKUKTKSKTKSNKOKNKMKLKKNKIKHKGKFKENKCNKAK@K?K>K=K<NK:K9K8K7K6K5K4K3K2K1K0K/K.NK,K+K*K)K(K'K&K%K$K#K"K!K KKKNKKKKKKNe]�(NKVKUNKSKRKSNKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?NK=K<K;K:K9K8NNK5K4K3K2K1K0K/K.K-K,NK*K)K(K'K&K%K$K#K"K!K KKKNKKKKKKKNe]�(NKUKTKSKRKQNKOKNKMKLKKKLNKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKNKKKKNe]�(NKTKSKRKQKPKOKNKMNKKKJNKHNKFKEKDKCKBKAK@K?NK=K<K;K:K9K8K7K6K5NK3K2K1K0K/K.K-K,K+K*K)K(K'NNK$K#K"K!K KKKKKKKKKKKKKNe]�(NKSKRKQKPKOKNKMKLKKKJKINKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"K!K KKKKKKKKKKKKKKNe]�(NKRKQKPKOKNKMKLKKKJKIKHKGKFNKDKCKBKAK@NK>K=K<K;K:K9K8K7NNK4K3NK1K0K/K.K-K,K+K*K)K(K'K&K%K$NK"K!K KKKKKKNKKKKKKKKNe]�(NKQKPKOKNKMNKMNKIKHKGKFKEKDKCKBKAK@K?K>NK<K;K:NK8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K KKKKKKKNKKKKKKKKNe]�(NKPKONKMKLKKKLKKKJKINKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!NKKKKKKKKKNKKKKKKKNe]�(NKOKNKMKLKKKJKKKLKKKJNKDKCKBKAKBNK>K=K<K;K:NK8NK6NK4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKNe]�(NKNKMKLKKKJKIKJKKNNKDNKBKAK@NK>K=K<K;K:K9NK7K6K5K4NK2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKNe]�(NKMKLKKKJKIKHNNKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5NK3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKNe]�(NKLKKKJNKHKGKFKEKDNKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKNe]�(NKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/NK-K,NK*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKNe]�(NKLKKKJKINKGKFNKDKCKBKAK@K?K>K=K<K;K:NK6K5K4K3K2NK0K/K.NK,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKNe]�(NKMNKKKJKINKGKFKEKDNKBKAK@K?K>K=K<K;NK5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKK
Ne]�(NKLKKKJKIKHKGKFKEKDNKBKAK@K?K>K=K<K;K:NK6K5K4K3NK1K0NK,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKKKK
K	Ne]�(NKKKJKIKHKGKFKEKDKCKBNK@NNK=K<K;K:K9K8K7K6NK2K1K0K/K.K-K,K+K*K)NNNNNNNNNNNNNNNNKKKKKKKKNKKKNKK
K	KNe]�(NKJKIKHKGKFNKDKCKBKAK@K?K>K=K<K;NK9K8K7K6K5NK3K2K1K0K/K.K-K,K+K*NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NKKKKKKKKKNKK
K	K
K	KKNe]�(NKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4NK2K1K0K/K.K-K,K+K*K)NK+K,K-K.K/K0K1K2K3K4K5K6K7K8NKKKKKKKKKKK
K	KK	KKKNe]�(NKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NK8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K)K*K+K,K-K.K/K0K1K2K3K4K5K6K7NKKKKKKKKKK
K	KKKKKKNe]�(NKIKHKGKFKENNNKAK@K?NK=NK;K:NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'NK+K,K-K.K/K0K1K2K3K4K5K6K7K8NKKKKKKKKNK	KKKKKKKNe]�(NKHKGKFKEKDKCNKAK@K?K>K=K<K;K:K9K8K7NK3K2K1K0K/K.K-K,K+K*K)K(K'K&NK,K-K.K/K0K1K2K3K4K5K6K7K8K9NKKKKKKKK
K	KKKKKKKKNe]�(NKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2NK.K-K,K+K*K)K(K'K&K%NK-K.K/K0K1K2K3K4K5K6K7K8K9K:NKKKKKKK
K	KKKKKKNKKNe]�(NKFNKDKCNKAK@K?NK=K<K;K:K9K8K7K6K5K4K3K2K1K0NK,K+K*K)K(K'K&K%K$NNNNNNNNNNNNNNNNKKKKKKKK
NKKKKNKK KNe]�(NKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK$K#K"K!K KKKKKKKKKKKKKKNNKKKKKNKKKKKK KK Ne]�(NKFNKDNKBKAK@K?K>NK<K;K:K9K8NK4K3K2K1K0K/K.K-K,NK*NK(NK&K%K$K#K"K!K KKKKKKKKKKKKKKKKKNKKNKKKKKKK KNe]�(NKGKFKEKDKCNKAK@K?NK;K:K9K8K7K6K5K4K3K2NK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKKKNKKKKKNKKNe]�(NKHNNKCKBNK@K?K>K=K<NK8K7K6K5K4K3K2K1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKNKK
K	KKKKKKKKNe]�(NKGKFKENKAK@K?K>K=K<K;K:K9K8K7K6K5NNK2NK0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K KKKKKKKKKKKNKKKKKKKNK	KNNKKKKNe]�(NKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK7K6K5K4NNK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKKNKK
K	KKKKKKNe]�(NKGKFKEKDKCKBKAK@K?NK=K<K;K:K9K8NK4K3K2K1K0NK.K-K,K+K*K)NK'K&K%K$K#K"K!K KKKKKKKKKKKKNKKKKKKKKK
K	KKKKKNe]�(NKHKGKFKEKDNKBKAK@K?K>NK:K9K8K7K6K5K4K3K2K1K0K/K.K-NK+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKNKKKKKKKKKNK	KKKKNe]�(NKIKHNKDKCKBKAK@K?K>K=K<K;NK9K8NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(NK&K%K$K#K"NK NKKKKKKKKKKKKKKKKKKKKK
K	KKKNe]�(NKHKGKFKEKDKCNKANK?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#NK!K KKKKNKKNKKKKKKKKKKKKKK
K	KK	Ne]�(NKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK8K7K6K5K4K3NK1K0K/NK-K,K+K*K)K(K'K&K%K$K#K"K!NKKKKKKKKKNKKKKNKKKKKKK
K	K
Ne]�(NKJKIKHKGKFKEKDKCKBKAK@K?K>K=NK;K:K9NK7K6K5NK3K2K1K0K1NK-K,K+K*K)NNK&NK$K#K"K!K KKKKKKKKKKKKKKKKKKKKKK
KNe]�(NKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:NK8K7K6NK4K3K2K1K0K/K.NK,K+K*K)K(K'K(NK$K#K"K!K KKKNKKKKKNKKNKKKKKKKKKNe]�(NKLKKKJKIKHKGKFKENKCKBKAK@NNNNK;K:K9K8K7K6K5NK3K2K1K0K/K.K-K,K+K*K)K(K)NK%K$K#K"K!K KKKKKNKKKKKKKKKKKKKKKNe]�(NKMKLKKKJKIKHNKFNKDKCKBKAK@K?K>K=K<K;K:NK8K7K6K7NK3K2K1NK/K.K-K,K+K*K)K(K'K&K%K$K#K"NK KKNKKNKKKNKKKKKKKKKKNe]�(NKNKMKLKKNKINKGKFKEKDKCKBKAK@K?K>K=NK;K:K9K8K7K6K5K4K3K2NK0K/K.K-K,K+K*K)K(K'K&K%NK#K"K!K KKKKKKKKNKKKKKKKKKKNe]�(NKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5NK3K2K1NK/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKKKNe]�(NKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%NK#K"K!K KKKKKKKKKKKKKKKKKNe]�(NKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8NK6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKNe]�(NKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKNe]�(NKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)NK'K&K%K$K#K"K!K KKKKKKKKKKKKKKNe]�(NKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;NK9K8NK6K5K4K3K2K1K0K/K.K-K,K+K*NK(K'NK%K$K#K"K!K KKKKKKKKKKKKKNe]�(NKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6NK4K3K2K1K0K/K.K-K,NK*K)K(NK&K%K$K#K"K!K KKKKKKKKKKKKNe]�(NKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*NK(K'K&K%K$K#K"K!K KKKKKKKKKKKNe]�(NKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7NNNNNNNNK.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKKKKKKKKNe]�(NKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8NK>K?K@KAKBKCNK/K.K-K,K+K*K)K(NK&K%NK#K"K!K KKKKKKKKKNe]�(NKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9NK=K>K?K@KAKBNK0K/K.K-K,K+K*K)K(K'K&NK$K#K"K!K KKKKKKKKNe]�(NKZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K;K<K=K>K?K@KANK1K0K/K.K-K,K+K*K)K(K'K(NK$K#NK!K KKKKKKKNe]�(NK[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;NK=K>K?K@KAKBNK2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K!K KKKKKKNe]�(NK\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<NK>K?K@KAKBKCNK3K2K1K0K/K.K-K,K+K*K)K(K'NK%K$K#K"K!K KKKKKNe]�(NK]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=NK?K@KAKBKCKDNK4K3K2K1K0K/K.K-K,K+NK)K(K'K&K%K$K#K"K!K KKKKNe]�(NK^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K?NNNNNNNK5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKKNe]�(NK_K^K]K\K[KZKYKXKWKVKUKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@K?K>K=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KK Ne]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej��  Kubaj�8  j[�  j��  M�Mj��  K ubj�9  j[�  j�9  Kj�9  �0.1.0�j�9  j�9  )��KYKE]�(K K K K ��K K K ����KKK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KLK�K�K���K K K ����KEK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KRK�K�K���K K K ����KPK�K�K���K K K ����KAK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KWK�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KGK�K�K���K K K ����KPK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KxK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KaK�K�K���K K K ����KoK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KlK�K�K���K K K ����KFK�K�K���K K K ����K K K K ��K K K ����KvK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KnK�K�K���K K K ����KwK�K�K���K K K ����KmK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KyK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KwK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K0K�K�K���K K K ����K K K K ��K K K ����KhK�K�K���K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K:K�K�K���K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KSK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KPK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K1K�K�K���K K K ����K2K�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����KRK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K9K�K�K���K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KBK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KFK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KKK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K|K�K��      K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.KdKdKd��K K K ����KTKdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K@KKYK���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����KTKKnK��K K K ����KSK�K�K���K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����K KdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKdKdKd��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����KTKKnK��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ������8      K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e��bj��  K,ub.