��      �Player�h ��)��}�(�level�K�exp�K#�recalcTimer�K �skills�}�(�3��	Abilities��Fireball����4�h
�Lightning_Bolt����7�h
�Ready_for_Battle����5�h
�Block����6�h
�Rending_Blow����1�h
�Charge����2�h
�Shocking_Grasp���u�
prevTarget�N�power�K�playerControlled���helmet��Items.Armors��Leather_Helm���)��}�(�armorVal�K
hK�
equippable���
consumable���weight�K�type�h"�color�]�(K�K�K�e�char��?��	throwable���name��Leather Helm�ub�armorPen�K �gold�KC�
healthTemp�K �dodge�K �	sightDist�K�
initiative�K�armor�h#�Cloth_Shirt���)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�Cloth Shirt�ub�leftHand��Items.Weapons��Tome���)��}�(hKh/h0h,�0H�h)�h*��addPower���range�Kh K h+K�magPower�K�
usesArrows��h-h.h4K h1�h2hBub�canMove���
countering���items�]�(�Items.Consumables��	GreenHerb���)��}�(h)�h*��healNum�Kh,h*h-h.h/�+�h2�
Green Herb�ubhQ)��}�(h)�h*�hTKh,h*h-h.h/hUh2hVubh%)��}�(h(K
hKh)�h*�h+K�pObject�Nh,h"h-h.h/h0h1�h2h3ubh#�	Iron_Helm���)��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�	Iron Helm�ubhA�Wooden_Shield���)��}�(hKh/h0h,�1H�h)�h*�hG�h(Kh K h+KhIK h-h.hHKhJ�h1�h2�Wooden Shield�ubh])��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2h`ubh])��}�(h(KhKh)�h*�h+Kh[Nh,h"h-h.h/h0h1�h2h`ubhA�	Longsword���)��}�(hKh/h0h,heh)�h*�hG�h[NhHKh Kh+KhIKhJ�h-h.h4Kh1�h2hkubhl)��}�(hKh/h0h,heh)�h*�hG�h[NhHKh Kh+KhIKhJ�h-h.h4Kh1�h2hkubhO�Scroll_of_Lightning_Bolt���)��}�(hKh)�h*��spell�hh[Nh,�scroll�h-h.h/�s�h2�Scroll of Lightning Bolt�ubhQ)��}�(h)�h*�hTKh[Nh,h*h-h.h/hUh2hVubh])��}�(h(KhKh)�h*�h+Kh[Nh,h"h-h.h/h0h1�h2h`ubhl)��}�(hKh/h0h,heh)�h*�hG�h[NhHKh Kh+KhIKhJ�h-h.h4Kh1�h2hkubh])��}�(h(KhKh)�h*�h+Kh[Nh,h"h-h.h/h0h1�h2h`ubh])��}�(h(KhKh)�h*�h+Kh[Nh,h"h-h.h/h0h1�h2h`ubhl)��}�(hKh/h0h,heh)�h*�hG�h[NhHKh Kh+KhIKhJ�h-h.h4Kh1�h2hkubhl)��}�(hKh/h0h,heh)�h*�hG�h[NhHKh Kh+KhIKhJ�h-h.h4Kh1�h2hkubhO�	Time_Bomb���)��}�(hKh/�o�h,h*h)�h*�h[N�dur�Kh-h.hHK h2�Bomb��desc��Explodes up after 3 turns��damage�K�radius�KubhA�Buckler���)��}�(hKh/h0h,hFh)�h*�hG�h(Kh K h+KhIK h-h.hHKhJ�h1�h2h�ubh])��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2h`ubhQ)��}�(h)�h*�hTKh,h*h-h.h/hUh2hVubh#�Chain_Shirt���)��}�(h(K#hKh)�h*�h+K#h,h:h-h.h/h0h1�h2�Chain Shirt�ubhl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4Kh1�h2hkubh])��}�(h(KhKh)�h*�h+Kh[Nh,h"h-h.h/h0h1�h2�+1 Iron Helm�ubh%)��}�(h(KhKh)�h*�h+Kh[Nh,h"h-h.h/h0h1�h2�+1 Leather Helm�ubhl)��}�(hKh/h0h,heh)�h*�hG�h[NhHKh Kh+KhIKhJ�h-h.h4K
h1�h2hkubhl)��}�(hKh/h0h,heh)�h*�hG�h[NhHKh Kh+KhIKhJ�h-h.h4K
h1�h2hkubh�)��}�(hKh/h�h,h*h)�h*�h[Nh�Kh-h.hHK h2h�h�h�h�Kh�Kubh])��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Iron Helm�ubhr)��}�(hKh)�h*�huhh,hvh-h.h/hwh2hxubhQ)��}�(h)�h*�hTK h,h*h-h.h/hUh2hVube�health�Kʌvisible���
baseHealth�M�	rightRing�N�accuracy�K �necklace�N�	rightHand�hA�
Greatsword���)��}�(hKh/h0h,�2H�h)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4Kh1�h2h�ubh/�@�h(K �
leftScroll�N�blocking���arrows�K�Class��Player_Classes��
Spellsword����	healthMax�M�leftRing�N�	recalcMax�K �healthCurve�G?�333333�rightScroll�N�invertColor���
hitEffects�]��skillLevels�}�(h	K hK hK hK hK hK hK uh[�Object�hғ�)��}�(�pLevel��LevelTypes.LevelTypes��Crypt���)��}�(�cLevel�K�args�]�(KKKKKKe�itemList�]�(hQhO�Bundle_Of_Arrows���h�hO�Scroll_of_Fireball���hrhA�Staff���hA�Iron_Shield���h�hbhlh�hA�Bow���hA�Spear���hA�Dagger���h<h#�	Cloth_Hat���h#�Leather_Shirt���h%h#�Iron_Breastplate���h]h�h#�
Chain_Helm���e�healingList�]�hQa�	equipList�]�(h�h�h�hbhlh�h�h�h�h<h�h�h%h�h]h�h�e�stairsUp�]�(K/K/e�	eliteList�]��Enemies.Undead��Cultist���a�Objects�}�(K@h�)��}�(h�h�h/h0�ID�K@�row�K>�col�K
h�hb)��}�(hKh/h0h,heh)�h*�hG�h[j  h(Kh K h+KhIK h-h.hHKhJ�h1�h2hfubh2�Item�ubKCh�)��}�(h�h�h/�x�j  KCj  K?j  K	h�h��Zombie���)��}�(hKhK h/j  �
dropChance�K(�
alliesList�]�(j  h�)��}�(h�h�h/j  j  KDj  K@j  K
h�j  )��}�(hKhK h/j  j  K(j  ]�(j  j  h�)��}�(h�h�h/j  j  KFj  KBj  K
h�j  )��}�(hKhK h/j  j  K(j  ]�(j  j  j  eh Kh!�h"h%)��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Leather Helm�ubh4K h5Kh6K h7K h8K	h9Kh�Kh@N�	cowardice�G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�+1 Leather Shirt�ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4K
h1�h2hkub�lastPlayerLoc�Nh(K �isAfraid��hh�K �lastPlayerMap�Nh�K�hearingDist�Kh�Nh͉h�]�h[j  �expNext�Kd�effects�]��
stealthVal�K h-]�(K�KKeh2j  ubh2�Enemy�ubeh Kh!�h"h%)��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Leather Helm�ubh4K h5K
h6K h7K h8K	h9Kh�Kh@Nj#  G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�+1 Leather Shirt�ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4K
h1�h2hkubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j  j/  Kdj0  ]�j2  K h-j3  h2j  ubh2j4  ubj  eh Kh!�h"h%)��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Leather Helm�ubh4K h5Kh6K h7K h8K	h9Kh�Kh@Nj#  G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�+1 Leather Shirt�ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4K
h1�h2hkubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j  j/  Kdj0  ]�j2  K h-j3  h2j  ubh2j4  ubKDj  KEh�)��}�(h�h�h/�=�j  KEj  KAj  K2hҌFeatures.Features��Chest���)��}�(hM]�h[jK  h-h.h/jM  h2jO  ubh2jO  ubKFj  KGh�)��}�(h�h�h/jM  j  KGj  KCj  K
h�jP  )��}�(hM]�(h�)��}�(hKh/h0h,h�h)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4K
h1�h2h�ubh�)��}�(h(KhKh)�h*�h+K
h,h"h-h.h/h0h1�h2�+1 Chain Helm�ubh�)��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Cloth Hat�ubhO�
Gold_Coins���)��}�(h)�h*�h,h*h-]�(K�K�Keh/�$��coins�Kh2�
Gold Coins�ubeh[jT  h-]�(KQKOKeh/jM  h2jO  ubh2jO  ubKHh�)��}�(h�h�h/�*�j  KHj  KDj  K,hҌLevelTypes.Decorations��Altar���)��}�(h2jn  h[jj  h/jl  ubh2jn  ubKIh�)��}�(h�h�h/h0j  KIj  K<j  K+h�h�h2h�ubKJh�)��}�(h�h�h/h0j  KJj  K<j  K+h�h�h2hkubKKh�)��}�(h�h�h/h�j  KKj  K<j  K+h�h�h2h�ubKLh�)��}�(h�h�h/h0j  KLj  K<j  K,h�h�h2h�ubKMh�)��}�(h�h�h/h0j  KMj  K<j  K,h�h�h2hkubK%h�)��}�(h�h�h/�E�j  K%j  Kj  KhҌFeatures.Stairs��	StairDown���)��}�(h�h�h[j|  j  J����j  K�moveCost�Kh�Nj  Kh2�Stairs�ubh2�Stairs Down�ubK&h�)��}�(h�h�h/jl  j  K&j  Kj  Kh�jm  �Ritual_Circle���)��}�(h2�Ritual Circle�h[j�  h/jl  ubh2j�  ubK'h�)��}�(h�h�h/j  j  K'j  Kj  Kh�h��Skeleton_Knight���)��}�(hKhK h/j  j  K(j  ]�(j�  h�)��}�(h�h�h/j  j  K(j  Kj  Kh�j�  )��}�(hKhK h/j  j  K(j  ]�(j�  j�  h�)��}�(h�h�h/�X�j  K)j  Kj  Kh�j  )��}�(hKhK h/j�  j  K(j  ]�(j�  j�  j�  eh Kh!�h"h�)��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Cloth Hat�ubh4K h5Kh6K h7K h8Kh9Kh�Kh@hC)��}�(hKh/h0h,hFh)�h*�hG�hHKh K h+KhIKhJ�h-h.h4K h1�h2hBubj#  G        hK�hL�hM]�h:h<)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�+1 Cloth Shirt�ubhHKh��h�Nh�K �cdMax�Kh�Nh�h�)��}�(hKh/h0h,h�h)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4K
h1�h2h�ubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j�  j/  Kdj0  ]�j2  K hTK h-j3  �cd�Kph2�Robed Cultist�ubh2j4  ubeh Kh!�h"h])��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Iron Helm�ubh4K h5Kh6K h7K h8Kh9Kh�Kh@hb)��}�(hKh/h0h,heh)�h*�hG�h(Kh K h+KhIK h-h.hHKhJ�h1�h2hfubj#  G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�+1 Leather Shirt�ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4K
h1�h2hkubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j�  j/  Kdj0  ]�j2  K h-j3  h2�Skeleton Knight�ubh2j4  ubj�  eh Kh!�h"h])��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Iron Helm�ubh4K h5Kh6K h7K h8Kh9Kh�Kh@hb)��}�(hKh/h0h,heh)�h*�hG�h(Kh K h+KhIK h-h.hHKhJ�h1�h2hfubj#  G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�+1 Leather Shirt�ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4K
h1�h2hkubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j�  j/  Kdj0  ]�j2  K h-j3  h2j�  ubh2j4  ubK(j�  K)j�  K*h�)��}�(h�h�h/j  j  K*j  Kj  K-h�j  )��}�(hKhK h/j  j  K(j  ]�j�  ah Kh!�h"h%)��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Leather Helm�ubh4K h5K	h6K h7K h8K	h9Kh�Kh@Nj#  G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�+1 Leather Shirt�ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4K
h1�h2hkubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j�  j/  Kdj0  ]�j2  K h-j3  h2j  ubh2j4  ubK+h�)��}�(h�h�h/j  j  K+j  Kj  Kh�j  )��}�(hKhK h/j  j  K(j  ]�(j�  h�)��}�(h�h�h/j  j  K4j  Kj  Kh�j�  )��}�(hKhK h/j  j  K(j  ]�(j�  j�  eh Kh!�h"h])��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Iron Helm�ubh4K h5Kh6K h7K h8Kh9Kh�Kh@hb)��}�(hKh/h0h,heh)�h*�hG�h(Kh K h+KhIK h-h.hHKhJ�h1�h2hfubj#  G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�+1 Leather Shirt�ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4K
h1�h2hkubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j�  j/  Kdj0  ]�j2  K h-j3  h2j�  ubh2j4  ubeh Kh!�h"h%)��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Leather Helm�ubh4K h5Kh6K h7K h8K	h9Kh�Kh@Nj#  G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�+1 Leather Shirt�ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4K
h1�h2hkubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j�  j/  Kdj0  ]�j2  K h-j3  h2j  ubh2j4  ubK,h�)��}�(h�h�h/jl  j  K,j  Kj  K,h�jo  )��}�(h2jn  h[j�  h/jl  ubh2jn  ubK-h�)��}�(h�h�h/jl  j  K-j  Kj  K-h�j�  )��}�(h2j�  h[j  h/jl  ubh2j�  ubK.h�)��}�(h�h�h/jl  j  K.j  Kj  K,h�jm  �Pile_of_Bones���)��}�(h2�Pile of Bones�h[j  h/jl  ubh2j  ubK/h�)��}�(h�h�h/jl  j  K/j  Kj  K-h�jo  )��}�(h2jn  h[j  h/jl  ubh2jn  ubK0h�)��}�(h�h�h/hUj  K0j  Kj  K
h�hQ)��}�(h)�h*�hTK h[j  h,h*h-h.h/hUh2hVubh2�Health�ubK1h�)��}�(h�h�h/jl  j  K1j  Kj  K,h�jo  )��}�(h2jn  h[j  h/jl  ubh2jn  ubK2h�)��}�(h�h�h/jl  j  K2j  Kj  K-h�j�  )��}�(h2j�  h[j  h/jl  ubh2j�  ubK3h�)��}�(h�h�h/j�  j  K3j  Kj  K1h�j  )��}�(hKhK h/j�  j  K(j  ]�j  ah Kh!�h"h�)��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Cloth Hat�ubh4K h5Kh6K h7K h8Kh9Kh�Kh@hC)��}�(hKh/h0h,hFh)�h*�hG�hHKh K h+KhIKhJ�h-h.h4K h1�h2hBubj#  G        hK�hL�hM]�h:h<)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�+1 Cloth Shirt�ubhHKh��h�Nh�K j�  Kh�Nh�h�)��}�(hKh/h0h,h�h)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4K
h1�h2h�ubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j  j/  Kdj0  ]�j2  K hTK h-j3  j�  Kph2j�  ubh2j4  ubK4j�  K5h�)��}�(h�h�h/j  j  K5j  K&j  Kh�j  )��}�(hKhK h/j  j  K(j  ]�j/  ah Kh!�h"h%)��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2�+1 Leather Helm�ubh4K h5Kh6K h7K h8K	h9Kh�Kh@Nj#  G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�+1 Leather Shirt�ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4K
h1�h2hkubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j/  j/  Kdj0  ]�j2  K h-j3  h2j  ubh2j4  ubK6h�)��}�(h�h�h/�S�j  K6j  K/j  K/h�j  �StairUp���)��}�(h[j?  h�h�j�  Kj  J����j  K/j  K/h�Nh2j�  ubh2�	Stairs Up�ubK7h�K8h�)��}�(h�h�h/jl  j  K8j  K0j  K*h�j�  )��}�(h2j�  h[jG  h/jl  ubh2j�  ubK9h�)��}�(h�h�h/�~�j  K9j  K4j  Kh�jN  �Brush���)��}�(h[jK  h-]�(KKnKeh/jM  h2jN  ubh2jN  ubK:h�)��}�(h�h�h/jM  j  K:j  K5j  K	h�jO  )��}�(h[jS  h-jR  h/jM  h2jN  ubh2jN  ubK;h�)��}�(h�h�h/jM  j  K;j  K5j  K
h�jO  )��}�(h[jW  h-jR  h/jM  h2jN  ubh2jN  ubK<h�)��}�(h�h�h/jM  j  K<j  K5j  Kh�jO  )��}�(h[j[  h-jR  h/jM  h2jN  ubh2jN  ubK=h�)��}�(h�h�h/jM  j  K=j  K5j  Kh�jO  )��}�(h[j_  h-jR  h/jM  h2jN  ubh2jN  ubK>h�)��}�(h�h�h/jM  j  K>j  K6j  K	h�jO  )��}�(h[jc  h-jR  h/jM  h2jN  ubh2jN  ubK?h�)��}�(h�h�h/hUj  K?j  K=j  K	h�hQ)��}�(h)�h*�hTK h[jg  h,h*h-h.h/hUh2hVubh2j  ubu�CollisionMap�]�(]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKK KKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKK KKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK K K KKKKKKKKKKKKKK KKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK K K KKKKKKKKKKKKKK KKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK KKKKKKKKKKKKKKKK KKKKKKKKKKKKKK KKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK KKKKKKKKKKKKKKKK KKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK KKKKKKKKKKKKKKKK KKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK KKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKK K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKK K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKee�djikstra_Stairs_Down�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKKK KKKKKKKKK	K
KKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKKKKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNK0K1K2K3K4K5K6NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNK/K0K1K2K3K4K5NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK	KKKKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNK.K/K0K1K2K3K4NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK
K	KKKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNK-K.K/K0K1K2K3NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK-K.K/K0K1K2K3NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK.K/K0K1K2K3K4NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK5NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK6NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK7NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK:K9K8NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK;NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK<NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK=NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKkKjKiKhKgKfKeNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKjKiKhKgKfKeKdKcKbKaK`K_K^K]K\K[KZKYKXKWKVKUNNNNNNNNNNNNNNNKCKBKAK@K?K@KAKBNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKkKjKiKhKgKfKeNNNNNNNNNNNNNNKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@KAKBKCNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKlKkKjKiKhKgKfNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKEKDKCKBKAKBKCKDNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKmKlKkKjKiKhKgNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKEKDKCKBKCKDKENNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKnKmKlKkKjKiKhNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKFKEKDKCKDKEKFNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKoKnKmKlKkKjKiNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKGKFKEKDKEKFKGNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKpKoKnKmKlKkKjNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKIKHKGKFKEKFKGKHNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKqKpKoKnKmKlKkNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKJKIKHKGKFKGKHKINNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKJKIKHKGKHKIKJNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�Tiles�}�(K }�(K �Tile�j  ��)��}�(h�h�j  ]�j  K j  K ubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubK	j  )��}�(h�h�j  ]�j  K j  K	ubK
j  )��}�(h�h�j  ]�j  K j  K
ubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubK j  )��}�(h�h�j  ]�j  K j  K ubK!j  )��}�(h�h�j  ]�j  K j  K!ubK"j  )��}�(h�h�j  ]�j  K j  K"ubK#j  )��}�(h�h�j  ]�j  K j  K#ubK$j  )��}�(h�h�j  ]�j  K j  K$ubK%j  )��}�(h�h�j  ]�j  K j  K%ubK&j  )��}�(h�h�j  ]�j  K j  K&ubK'j  )��}�(h�h�j  ]�j  K j  K'ubK(j  )��}�(h�h�j  ]�j  K j  K(ubK)j  )��}�(h�h�j  ]�j  K j  K)ubK*j  )��}�(h�h�j  ]�j  K j  K*ubK+j  )��}�(h�h�j  ]�j  K j  K+ubK,j  )��}�(h�h�j  ]�j  K j  K,ubK-j  )��}�(h�h�j  ]�j  K j  K-ubK.j  )��}�(h�h�j  ]�j  K j  K.ubK/j  )��}�(h�h�j  ]�j  K j  K/ubK0j  )��}�(h�h�j  ]�j  K j  K0ubK1j  )��}�(h�h�j  ]�j  K j  K1ubK2j  )��}�(h�h�j  ]�j  K j  K2ubK3j  )��}�(h�h�j  ]�j  K j  K3ubK4j  )��}�(h�h�j  ]�j  K j  K4ubK5j  )��}�(h�h�j  ]�j  K j  K5ubK6j  )��}�(h�h�j  ]�j  K j  K6ubK7j  )��}�(h�h�j  ]�j  K j  K7ubK8j  )��}�(h�h�j  ]�j  K j  K8ubK9j  )��}�(h�h�j  ]�j  K j  K9ubK:j  )��}�(h�h�j  ]�j  K j  K:ubK;j  )��}�(h�h�j  ]�j  K j  K;ubK<j  )��}�(h�h�j  ]�j  K j  K<ubK=j  )��}�(h�h�j  ]�j  K j  K=ubK>j  )��}�(h�h�j  ]�j  K j  K>ubK?j  )��}�(h�h�j  ]�j  K j  K?ubK@j  )��}�(h�h�j  ]�j  K j  K@ubKAj  )��}�(h�h�j  ]�j  K j  KAubKBj  )��}�(h�h�j  ]�j  K j  KBubKCj  )��}�(h�h�j  ]�j  K j  KCubKDj  )��}�(h�h�j  ]�j  K j  KDubKEj  )��}�(h�h�j  ]�j  K j  KEubKFj  )��}�(h�h�j  ]�j  K j  KFubKGj  )��}�(h�h�j  ]�j  K j  KGubKHj  )��}�(h�h�j  ]�j  K j  KHubKIj  )��}�(h�h�j  ]�j  K j  KIubKJj  )��}�(h�h�j  ]�j  K j  KJubKKj  )��}�(h�h�j  ]�j  K j  KKubKLj  )��}�(h�h�j  ]�j  K j  KLubKMj  )��}�(h�h�j  ]�j  K j  KMubKNj  )��}�(h�h�j  ]�j  K j  KNubKOj  )��}�(h�h�j  ]�j  K j  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�K%aj  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�K&aj  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�K'aj  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�K(aj  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�K)aj  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK	}�(K j  )��}�(h�h�j  ]�j  K	j  K ubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubK	j  )��}�(h�h�j  ]�j  K	j  K	ubK
j  )��}�(h�h�j  ]�j  K	j  K
ubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubKj  )��}�(h�h�j  ]�j  K	j  KubK j  )��}�(h�h�j  ]�j  K	j  K ubK!j  )��}�(h�h�j  ]�j  K	j  K!ubK"j  )��}�(h�h�j  ]�j  K	j  K"ubK#j  )��}�(h�h�j  ]�j  K	j  K#ubK$j  )��}�(h�h�j  ]�j  K	j  K$ubK%j  )��}�(h�h�j  ]�j  K	j  K%ubK&j  )��}�(h�h�j  ]�j  K	j  K&ubK'j  )��}�(h�h�j  ]�j  K	j  K'ubK(j  )��}�(h�h�j  ]�j  K	j  K(ubK)j  )��}�(h�h�j  ]�j  K	j  K)ubK*j  )��}�(h�h�j  ]�j  K	j  K*ubK+j  )��}�(h�h�j  ]�j  K	j  K+ubK,j  )��}�(h�h�j  ]�j  K	j  K,ubK-j  )��}�(h�h�j  ]�j  K	j  K-ubK.j  )��}�(h�h�j  ]�j  K	j  K.ubK/j  )��}�(h�h�j  ]�j  K	j  K/ubK0j  )��}�(h�h�j  ]�j  K	j  K0ubK1j  )��}�(h�h�j  ]�j  K	j  K1ubK2j  )��}�(h�h�j  ]�j  K	j  K2ubK3j  )��}�(h�h�j  ]�j  K	j  K3ubK4j  )��}�(h�h�j  ]�j  K	j  K4ubK5j  )��}�(h�h�j  ]�j  K	j  K5ubK6j  )��}�(h�h�j  ]�j  K	j  K6ubK7j  )��}�(h�h�j  ]�j  K	j  K7ubK8j  )��}�(h�h�j  ]�j  K	j  K8ubK9j  )��}�(h�h�j  ]�j  K	j  K9ubK:j  )��}�(h�h�j  ]�j  K	j  K:ubK;j  )��}�(h�h�j  ]�j  K	j  K;ubK<j  )��}�(h�h�j  ]�j  K	j  K<ubK=j  )��}�(h�h�j  ]�j  K	j  K=ubK>j  )��}�(h�h�j  ]�j  K	j  K>ubK?j  )��}�(h�h�j  ]�j  K	j  K?ubK@j  )��}�(h�h�j  ]�j  K	j  K@ubKAj  )��}�(h�h�j  ]�j  K	j  KAubKBj  )��}�(h�h�j  ]�j  K	j  KBubKCj  )��}�(h�h�j  ]�j  K	j  KCubKDj  )��}�(h�h�j  ]�j  K	j  KDubKEj  )��}�(h�h�j  ]�j  K	j  KEubKFj  )��}�(h�h�j  ]�j  K	j  KFubKGj  )��}�(h�h�j  ]�j  K	j  KGubKHj  )��}�(h�h�j  ]�j  K	j  KHubKIj  )��}�(h�h�j  ]�j  K	j  KIubKJj  )��}�(h�h�j  ]�j  K	j  KJubKKj  )��}�(h�h�j  ]�j  K	j  KKubKLj  )��}�(h�h�j  ]�j  K	j  KLubKMj  )��}�(h�h�j  ]�j  K	j  KMubKNj  )��}�(h�h�j  ]�j  K	j  KNubKOj  )��}�(h�h�j  ]�j  K	j  KOubuK
}�(K j  )��}�(h�h�j  ]�j  K
j  K ubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubK	j  )��}�(h�h�j  ]�j  K
j  K	ubK
j  )��}�(h�h�j  ]�j  K
j  K
ubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  �      K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubKj  )��}�(h�h�j  ]�j  K
j  KubK j  )��}�(h�h�j  ]�j  K
j  K ubK!j  )��}�(h�h�j  ]�j  K
j  K!ubK"j  )��}�(h�h�j  ]�j  K
j  K"ubK#j  )��}�(h�h�j  ]�j  K
j  K#ubK$j  )��}�(h�h�j  ]�j  K
j  K$ubK%j  )��}�(h�h�j  ]�j  K
j  K%ubK&j  )��}�(h�h�j  ]�j  K
j  K&ubK'j  )��}�(h�h�j  ]�j  K
j  K'ubK(j  )��}�(h�h�j  ]�j  K
j  K(ubK)j  )��}�(h�h�j  ]�j  K
j  K)ubK*j  )��}�(h�h�j  ]�j  K
j  K*ubK+j  )��}�(h�h�j  ]�j  K
j  K+ubK,j  )��}�(h�h�j  ]�j  K
j  K,ubK-j  )��}�(h�h�j  ]�j  K
j  K-ubK.j  )��}�(h�h�j  ]�j  K
j  K.ubK/j  )��}�(h�h�j  ]�j  K
j  K/ubK0j  )��}�(h�h�j  ]�j  K
j  K0ubK1j  )��}�(h�h�j  ]�j  K
j  K1ubK2j  )��}�(h�h�j  ]�j  K
j  K2ubK3j  )��}�(h�h�j  ]�j  K
j  K3ubK4j  )��}�(h�h�j  ]�j  K
j  K4ubK5j  )��}�(h�h�j  ]�j  K
j  K5ubK6j  )��}�(h�h�j  ]�j  K
j  K6ubK7j  )��}�(h�h�j  ]�j  K
j  K7ubK8j  )��}�(h�h�j  ]�j  K
j  K8ubK9j  )��}�(h�h�j  ]�j  K
j  K9ubK:j  )��}�(h�h�j  ]�j  K
j  K:ubK;j  )��}�(h�h�j  ]�j  K
j  K;ubK<j  )��}�(h�h�j  ]�j  K
j  K<ubK=j  )��}�(h�h�j  ]�j  K
j  K=ubK>j  )��}�(h�h�j  ]�j  K
j  K>ubK?j  )��}�(h�h�j  ]�j  K
j  K?ubK@j  )��}�(h�h�j  ]�j  K
j  K@ubKAj  )��}�(h�h�j  ]�j  K
j  KAubKBj  )��}�(h�h�j  ]�j  K
j  KBubKCj  )��}�(h�h�j  ]�j  K
j  KCubKDj  )��}�(h�h�j  ]�j  K
j  KDubKEj  )��}�(h�h�j  ]�j  K
j  KEubKFj  )��}�(h�h�j  ]�j  K
j  KFubKGj  )��}�(h�h�j  ]�j  K
j  KGubKHj  )��}�(h�h�j  ]�j  K
j  KHubKIj  )��}�(h�h�j  ]�j  K
j  KIubKJj  )��}�(h�h�j  ]�j  K
j  KJubKKj  )��}�(h�h�j  ]�j  K
j  KKubKLj  )��}�(h�h�j  ]�j  K
j  KLubKMj  )��}�(h�h�j  ]�j  K
j  KMubKNj  )��}�(h�h�j  ]�j  K
j  KNubKOj  )��}�(h�h�j  ]�j  K
j  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�K*aj  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�K+aj  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�K,aj  Kj  K,ubK-j  )��}�(h�h�j  ]�K-aj  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�K.aj  Kj  K,ubK-j  )��}�(h�h�j  ]�K/aj  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�K0aj  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�K1aj  Kj  K,ubK-j  )��}�(h�h�j  ]�K2aj  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�K3aj  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�K4aj  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(�      h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK}�(K j  )��}�(h�h�j  ]�j  Kj  K ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK	j  )��}�(h�h�j  ]�j  Kj  K	ubK
j  )��}�(h�h�j  ]�j  Kj  K
ubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubKj  )��}�(h�h�j  ]�j  Kj  KubK j  )��}�(h�h�j  ]�j  Kj  K ubK!j  )��}�(h�h�j  ]�j  Kj  K!ubK"j  )��}�(h�h�j  ]�j  Kj  K"ubK#j  )��}�(h�h�j  ]�j  Kj  K#ubK$j  )��}�(h�h�j  ]�j  Kj  K$ubK%j  )��}�(h�h�j  ]�j  Kj  K%ubK&j  )��}�(h�h�j  ]�j  Kj  K&ubK'j  )��}�(h�h�j  ]�j  Kj  K'ubK(j  )��}�(h�h�j  ]�j  Kj  K(ubK)j  )��}�(h�h�j  ]�j  Kj  K)ubK*j  )��}�(h�h�j  ]�j  Kj  K*ubK+j  )��}�(h�h�j  ]�j  Kj  K+ubK,j  )��}�(h�h�j  ]�j  Kj  K,ubK-j  )��}�(h�h�j  ]�j  Kj  K-ubK.j  )��}�(h�h�j  ]�j  Kj  K.ubK/j  )��}�(h�h�j  ]�j  Kj  K/ubK0j  )��}�(h�h�j  ]�j  Kj  K0ubK1j  )��}�(h�h�j  ]�j  Kj  K1ubK2j  )��}�(h�h�j  ]�j  Kj  K2ubK3j  )��}�(h�h�j  ]�j  Kj  K3ubK4j  )��}�(h�h�j  ]�j  Kj  K4ubK5j  )��}�(h�h�j  ]�j  Kj  K5ubK6j  )��}�(h�h�j  ]�j  Kj  K6ubK7j  )��}�(h�h�j  ]�j  Kj  K7ubK8j  )��}�(h�h�j  ]�j  Kj  K8ubK9j  )��}�(h�h�j  ]�j  Kj  K9ubK:j  )��}�(h�h�j  ]�j  Kj  K:ubK;j  )��}�(h�h�j  ]�j  Kj  K;ubK<j  )��}�(h�h�j  ]�j  Kj  K<ubK=j  )��}�(h�h�j  ]�j  Kj  K=ubK>j  )��}�(h�h�j  ]�j  Kj  K>ubK?j  )��}�(h�h�j  ]�j  Kj  K?ubK@j  )��}�(h�h�j  ]�j  Kj  K@ubKAj  )��}�(h�h�j  ]�j  Kj  KAubKBj  )��}�(h�h�j  ]�j  Kj  KBubKCj  )��}�(h�h�j  ]�j  Kj  KCubKDj  )��}�(h�h�j  ]�j  Kj  KDubKEj  )��}�(h�h�j  ]�j  Kj  KEubKFj  )��}�(h�h�j  ]�j  Kj  KFubKGj  )��}�(h�h�j  ]�j  Kj  KGubKHj  )��}�(h�h�j  ]�j  Kj  KHubKIj  )��}�(h�h�j  ]�j  Kj  KIubKJj  )��}�(h�h�j  ]�j  Kj  KJubKKj  )��}�(h�h�j  ]�j  Kj  KKubKLj  )��}�(h�h�j  ]�j  Kj  KLubKMj  )��}�(h�h�j  ]�j  Kj  KMubKNj  )��}�(h�h�j  ]�j  Kj  KNubKOj  )��}�(h�h�j  ]�j  Kj  KOubuK }�(K j  )��}�(h�h�j  ]�j  K j  K ubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubK	j  )��}�(h�h�j  ]�j  K j  K	ubK
j  )��}�(h�h�j  ]�j  K j  K
ubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubKj  )��}�(h�h�j  ]�j  K j  KubK j  )��}�(h�h�j  ]�j  K j  K ubK!j  )��}�(h�h�j  ]�j  K j  K!ubK"j  )��}�(h�h�j  ]�j  K j  K"ubK#j  )��}�(h�h�j  ]�j  K j  K#ubK$j  )��}�(h�h�j  ]�j  K j  K$ubK%j  )��}�(h�h�j  ]�j  K j  K%ubK&j  )��}�(h�h�j  ]�j  K j  K&ubK'j  )��}�(h�h�j  ]�j  K j  K'ubK(j  )��}�(h�h�j  ]�j  K j  K(ubK)j  )��}�(h�h�j  ]�j  K j  K)ubK*j  )��}�(h�h�j  ]�j  K j  K*ubK+j  )��}�(h�h�j  ]�j  K j  K+ubK,j  )��}�(h�h�j  ]�j  K j  K,ubK-j  )��}�(h�h�j  ]�j  K j  K-ubK.j  )��}�(h�h�j  ]�j  K j  K.ubK/j  )��}�(h�h�j  ]�j  K j  K/ubK0j  )��}�(h�h�j  ]�j  K j  K0ubK1j  )��}�(h�h�j  ]�j  K j  K1ubK2j  )��}�(h�h�j  ]�j  K j  K2ubK3j  )��}�(h�h�j  ]�j  K j  K3ubK4j  )��}�(h�h�j  ]�j  K j  K4ubK5j  )��}�(h�h�j  ]�j  K j  K5ubK6j  )��}�(h�h�j  ]�j  K j  K6ubK7j  )��}�(h�h�j  ]�j  K j  K7ubK8j  )��}�(h�h�j  ]�j  K j  K8ubK9j  )��}�(h�h�j  ]�j  K j  K9ubK:j  )��}�(h�h�j  ]�j  K j  K:ubK;j  )��}�(h�h�j  ]�j  K j  K;ubK<j  )��}�(h�h�j  ]�j  K j  K<ubK=j  )��}�(h�h�j  ]�j  K j  K=ubK>j  )��}�(h�h�j  ]�j  K j  K>ubK?j  )��}�(h�h�j  ]�j  K j  K?ubK@j  )��}�(h�h�j  ]�j  K j  K@ubKAj  )��}�(h�h�j  ]�j  K j  KAubKBj  )��}�(h�h�j  ]�j  K j  KBubKCj  )��}�(h�h�j  ]�j  K j  KCubKDj  )��}�(h�h�j  ]�j  K j  KDubKEj  )��}�(h�h�j  ]�j  K j  KEubKFj  )��}�(h�h�j  ]�j  K j  KFubKGj  )��}�(h�h�j  ]�j  K j  KGubKHj  )��}�(h�h�j  ]�j  K j  KHubKIj  )��}�(h�h�j  ]�j  K j  KIubKJj  )��}�(h�h�j  ]�j  K j  KJubKKj  )��}�(h�h�j  ]�j  K j  KKubKLj  )��}�(h�h�j  ]�j  K j  KLubKMj  )��}�(h�h�j  ]�j  K j  KMubKNj  )��}�(h�h�j  ]�j  K j  KNubKOj  )��}�(h�h�j  ]�j  K j  KOubuK!}�(K j  )��}�(h�h�j  ]�j  K!j  K ubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubK	j  )��}�(h�h�j  ]�j  K!j  K	ubK
j  )��}�(h�h�j  ]�j  K!j  K
ubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubKj  )��}�(h�h�j  ]�j  K!j  KubK j  )��}�(h�h�j  ]�j  K!j  K ubK!j  )��}�(h�h�j  ]�j  K!j  K!ubK"j  )��}�(h�h�j  ]�j  K!j  K"ubK#j  )��}�(h�h�j  ]�j  K!j  K#ubK$j  )��}�(h�h�j  ]�j  K!j  K$ubK%j  )��}�(h�h�j  ]�j  K!j  K%ubK&j  )��}�(h�h�j  ]�j  K!j  K&ubK'j  )��}�(h�h�j  ]�j  K!j  K'ubK(j  )��}�(h�h�j  ]�j  K!j  K(ubK)j  )��}�(h�h�j  ]�j  K!j  K)ubK*j  )��}�(h�h�j  ]�j  K!j  K*ubK+j  )��}�(h�h�j  ]�j  K!j  K+ubK,j  )��}�(h�h�j  ]�j  K!j  K,ubK-j  )��}�(h�h�j  ]�j  K!j  K-ubK.j  )��}�(h�h�j  ]�j  K!j  K.ubK/j  )��}�(h�h�j  ]�j  K!j  K/ubK0j  )��}�(h�h�j  ]�j  K!j  K0ubK1j  )��}�(h�h�j  ]�j  K!j  K1ubK2j  )��}�(h�h�j  ]�j  K!j  K2ubK3j  )��}�(h�h�j  ]�j  K!j  K3ubK4j  )��}�(h�h�j  ]�j  K!j  K4ubK5j  )��}�(h�h�j  ]�j  K!j  K5ubK6j  )��}�(h�h�j  ]�j  K!j  K6ubK7j  )��}�(h�h�j  ]�j  K!j  K7ubK8j  )��}�(h�h�j  ]�j  K!j  K8ubK9j  )��}�(h�h�j  ]�j  K!j  K9ubK:j  )��}�(h�h�j  ]�j  K!j  K:ubK;j  )��}�(h�h�j  ]�j  K!j  K;ubK<j  )��}�(h�h�j  ]�j  K!j  K<ubK=j  )��}�(h�h�j  ]�j  K!j  K=ubK>j  )��}�(h�h�j  ]�j  K!j  K>ubK?j  )��}�(h�h�j  ]�j  K!j  K?ubK@j  )��}�(h�h�j  ]�j  K!j  K@ubKAj  )��}�(h�h�j  ]�j  K!j  KAubKBj  )��}�(h�h�j  ]�j  K!j  KBubKCj  )��}�(h�h�j  ]�j  K!j  KCubKDj  )��}�(h�h�j  ]�j  K!j  KDubKEj  )��}�(h�h�j  ]�j  K!j  KEubKFj  )��}�(h�h�j  ]�j  K!j  KFubKGj  )��}�(h�h�j  ]�j  K!j  KGubKHj  )��}�(h�h�j  ]�j  K!j  KHubKIj  )��}�(h�h�j  ]�j  K!j  KIubKJj  )��}�(h�h�j  ]�j  K!j  KJubKKj  )��}�(h�h�j  ]�j  K!j  KKubKLj  )��}�(h�h�j  ]�j  K!j  KLubKMj  )��}�(h�h�j  ]�j  K!j  KMubKNj  )��}�(h�h�j  ]�j  K!j  KNubKOj  )��}�(h�h�j  ]�j  K!j  KOubuK"}�(K j  )��}�(h�h�j  ]�j  K"j  K ubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubK	j  )��}�(h�h�j  ]�j  K"j  K	ubK
j  )��}�(h�h�j  ]�j  K"j  K
ubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubKj  )��}�(h�h�j  ]�j  K"j  KubK j  )��}�(h�h�j  ]�j  K"j  K ubK!j  )��}�(h�h�j  ]�j  K"j  K!ubK"j  )��}�(h�h�j  ]�j  K"j  K"ubK#j  )��}�(h�h�j  ]�j  K"j  K#ubK$j  )��}�(h�h�j  ]�j  K"j  K$ubK%j  )��}�(h�h�j  ]�j  K"j  K%ubK&j  )��}�(h�h�j  ]�j  K"j  K&ubK'j  )��}�(h�h�j  ]�j  K"j  K'ubK(j  )��}�(h�h�j  ]�j  K"j  K(ubK)j  )��}�(h�h�j  ]�j  K"j  K)ubK*j  )��}�(h�h�j  ]�j  K"j  K*ubK+j  )��}�(h�h�j  ]�j  K"j  K+ubK,j  )��}�(h�h�j  ]�j  K"j  K,ubK-j  )��}�(h�h�j  ]�j  K"j  K-ubK.j  )��}�(h�h�j  ]�j  K"j  K.ubK/j  )��}�(h�h�j  ]�j  K"j  K/ubK0j  )��}�(h�h�j  ]�j  K"j  K0ubK1j  )��}�(h�h�j  ]�j  K"j  K1ubK2j  )��}�(h�h�j  ]�j  K"j  K2ubK3j  )��}�(h�h�j  ]�j  K"j  K3ubK4j  )��}�(h�h�j  ]�j  K"j  K4ubK5j  )��}�(h�h�j  ]�j  K"j  K5ubK6j  )��}�(h�h�j  ]�j  K"j  K6ubK7j  )��}�(h�h�j  ]�j  K"j  K7ubK8j  )��}�(h�h�j  ]�j  K"j  K8ubK9j  )��}�(h�h�j  ]�j  K"j  K9ubK:j  )��}�(h�h�j  ]�j  K"j  K:ubK;j  )��}�(h�h�j  ]�j  K"j  K;ubK<j  )��}�(h�h�j  ]�j  K"j  K<ubK=j  )��}�(h�h�j  ]�j  K"j  K=ubK>j  )��}�(h�h�j  ]�j  K"j  K>ubK?j  )��}�(h�h�j  ]�j  K"j  K?ubK@j  )��}�(h�h�j  ]�j  K"j  K@ubKAj  )��}�(h�h�j  ]�j  K"j  KAubKBj  )��}�(h�h�j  ]�j  K"j  KBubKCj  )��}�(h�h�j  ]�j  K"j  KCubKDj  )��}�(h�h�j  ]�j  K"j  KDubKEj  )��}�(h�h�j  ]�j  K"j  KEubKFj  )��}�(h�h�j  ]�j  K"j  KFubKGj  )��}�(h�h�j  ]�j  K"j  KGubKHj  )��}�(h�h�j  ]�j  K"j  KHubKIj  )��}�(h�h�j  ]�j  K"j  KIubKJj  )��}�(h�h�j  ]�j  K"j  KJubKKj  )��}�(h�h�j  ]�j  K"j  KKubKLj  )��}�(h�h�j  ]�j  K"j  KLubKMj  )��}�(h�h�j  ]�j  K"j  KMubKNj  )��}�(h�h�j  ]�j  K"j  KNubKOj  )��}�(h�h�j  ]�j  K"j  KOubuK#}�(K j  )��}�(h�h�j  ]�j  K#j  K ubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubK	j  )��}�(h�h�j  ]�j  K#j  K	ubK
j  )��}�(h�h�j  ]�j  K#j  K
ubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubKj  )��}�(h�h�j  ]�j  K#j  KubK j  )��}�(h�h�j  ]�j  K#j  K ubK!j  )��}�(h�h�j  ]�j  K#j  K!ubK"j  )��}�(h�h�j  ]�j  K#j  K"ubK#j  )��}�(h�h�j  ]�j  K#j  K#ubK$j  )��}�(h�h�j  ]�j  K#j  K$ubK%j  )��}�(h�h�j  ]�j  K#j  K%ubK&j  )��}�(h�h�j  ]�j  K#j  K&ubK'j  )��}�(h�h�j  ]�j  K#j  K'ubK(j  )��}�(h�h�j  ]�j  K#j  K(ubK)j  )��}�(h�h�j  ]�j  K#j  K)ubK*j  )��}�(h�h�j  ]�j  K#j  K*ubK+j  )��}�(h�h�j  ]�j  K#j  K+ubK,j  )��}�(h�h�j  ]�j  K#j  K,ubK-j  )��}�(h�h�j  ]�j  K#j  K-ubK.j  )��}�(h�h�j  ]�j  K#j  K.ubK/j  )��}�(h�h�j  ]�j  K#j  K/ubK0j  )��}�(h�h�j  ]�j  K#j  K0ubK1j  )��}�(h�h�j  ]�j  K#j  K1ubK2j  )��}�(h�h�j  ]�j  K#j  K2ubK3j  )��}�(h�h�j  ]�j  K#j  K3ubK4j  )��}�(h�h�j  ]�j  K#j  K4ubK5j  )��}�(h�h�j  ]�j  K#j  K5ubK6j  )��}�(h�h�j  ]�j  K#j  K6ubK7j  )��}�(h�h�j  ]�j  K#j  K7ubK8j  )��}�(h�h�j  ]�j  K#j  K8ubK9j  )��}�(h�h�j  ]�j  K#j  K9ubK:j  )��}�(h�h�j  ]�j  K#j  K:ubK;j  )��}�(h�h�j  ]�j  K#j  K;ubK<j  )��}�(h�h�j  ]�j  K#j  K<ubK=j  )��}�(h�h�j  ]�j  K#j  K=ubK>j  )��}�(h�h�j  ]�j  K#j  K>ubK?j  )��}�(h�h�j  ]�j  K#j  K?ubK@j  )��}�(h�h�j  ]�j  K#j  K@ubKAj  )��}�(h�h�j  ]�j  K#j  KAubKBj  )��}�(h�h�j  ]�j  K#j  KBubKCj  )��}�(h�h�j  ]�j  K#j  KCubKDj  )��}�(h�h�j  ]�j  K#j  KDubKEj  )��}�(h�h�j  ]�j  K#j  KEubKFj  )��}�(h�h�j  ]�j  K#j  KFubKGj  )��}�(h�h�j  ]�j  K#j  KGubKHj  )��}�(h�h�j  ]�j  K#j  KHubKIj  )��}�(h�h�j  ]�j  K#j  KIubKJj  )��}�(h�h�j  ]�j  K#j  KJubKKj  )��}�(h�h�j  ]�j  K#j  KKubKLj  )��}�(h�h�j  ]�j  K#j  KLubKMj  )��}�(h�h�j  ]�j  K#j  KMubKNj  )��}�(h�h�j  ]�j  K#j  KNubKOj  )��}�(h�h�j  ]�j  K#j  KOubuK$}�(K j  )��}�(h�h�j  ]�j  K$j  K ubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubK	j  )��}�(h�h�j  ]�j  K$j  K	ubK
j  )��}�(h�h�j  ]�j  K$j  K
ubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubKj  )��}�(h�h�j  ]�j  K$j  KubK j  )��}�(h�h�j  ]�j  K$j  K ubK!j  )��}�(h�h�j  ]�j  K$j  K!ubK"j  )��}�(h�h�j  ]�j  K$j  K"ubK#j  )��}�(h�h�j  ]�j  K$j  K#ubK$j  )��}�(h�h�j  ]�j  K$j  K$ubK%j  )��}�(h�h�j  ]�j  K$j  K%ubK&j  )��}�(h�h�j  ]�j  K$j  K&ubK'j  )��}�(h�h�j  ]�j  K$j  K'ubK(j  )��}�(h�h�j  ]�j  K$j  K(ubK)j  )��}�(h�h�j  ]�j  K$j  K)ubK*j  )��}�(h�h�j  ]�j  K$j  K*ubK+j  )��}�(h�h�j  ]�j  K$j  K+ubK,j  )��}�(h�h�j  ]�j  K$j  K,ubK-j  )��}�(h�h�j  ]�j  K$j  K-ubK.j  )��}�(h�h�j  ]�j  K$j  K.ubK/j  )��}�(h�h�j  ]�j  K$j  K/ubK0j  )��}�(h�h�j  ]�j  K$j  K0ubK1j  )��}�(h�h�j  ]�j  K$j  K1ubK2j  )��}�(h�h�j  ]�j  K$j  K2ubK3j  )��}�(h�h�j  ]�j  K$j  K3ubK4j  )��}�(h�h�j  ]�j  K$j  K4ubK5j  )��}�(h�h�j  ]�j  K$j  K5ubK6j  )��}�(h�h�j  ]�j  K$j  K6ubK7j  )��}�(h�h�j  ]�j  K$j  K7ubK8j  )��}�(h�h�j  ]�j  K$j  K8ubK9j  )��}�(h�h�j  ]�j  K$j  K9ubK:j  )��}�(h�h�j  ]�j  K$j  K:ubK;j  )��}�(h�h�j  ]�j  K$j  K;ubK<j  )��}�(h�h�j  ]�j  K$j  K<ubK=j  )��}�(h�h�j  ]�j  K$j  K=ubK>j  )��}�(h�h�j  ]�j  K$j  K>ubK?j  )��}�(h�h�j  ]�j  K$j  K?ubK@j  )��}�(h�h�j  ]�j  K$j  K@ubKAj  )��}�(h�h�j  ]�j  K$j  KAubKBj  )��}�(h�h�j  ]�j  K$j  KBubKCj  )��}�(h�h�j  ]�j  K$j  KCubKDj  )��}�(h�h�j  ]�j  K$j  KDubKEj  )��}�(h�h�j  ]�j  K$j  KEubKFj  )��}�(h�h�j  ]�j  K$j  KFubKGj  )��}�(h�h�j  ]�j  K$j  KGubKHj  )��}�(h�h�j  ]�j  K$j  KHubKIj  )��}�(h�h�j  ]�j  K$j  KIubKJj  )��}�(h�h�j  ]�j  K$j  KJubKKj  )��}�(h�h�j  ]�j  K$j  KKubKLj  )��}�(h�h�j  ]�j  K$j  KLubKMj  )��}�(h�h�j  ]�j  K$j  KMubKNj  )��}�(h�h�j  ]�j  K$j  KNubKOj  )��}�(h�h�j  ]�j  K$j  KOubuK%}�(K j  )��}�(h�h�j  ]�j  K%j  K ubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubK	j  )��}�(h�h�j  ]�j  K%j  K	ubK
j  )��}�(h�h�j  ]�j  K%j  K
ubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubKj  )��}�(h�h�j  ]�j  K%j  KubK j  )��}�(h�h�j  ]�j  K%j  K ubK!j  )��}�(h�h�j  ]�j  K%j  K!ubK"j  )��}�(h�h�j  ]�j  K%j  K"ubK#j  )��}�(h�h�j  ]�j  K%j  K#ubK$j  )��}�(h�h�j  ]�j  K%j  K$ubK%j  )��}�(h�h�j  ]�j  K%j  K%ubK&j  )��}�(h�h�j  ]�j  K%j  K&ubK'j  )��}�(h�h�j  ]�j  K%j  K'ubK(j  )��}�(h�h�j  ]�j  K%j  K(ubK)j  )��}�(h�h�j  ]�j  K%j  K)ubK*j  )��}�(h�h�j  ]�j  K%j  K*ubK+j  )��}�(h�h�j  ]�j  K%j  K+ubK,j  )��}�(h�h�j  ]�j  K%j  K,ubK-j  )��}�(h�h�j  ]�j  K%j  K-ubK.j  )��}�(h�h�j  ]�j  K%j  K.ubK/j  )��}�(h�h�j  ]�j  K%j  K/ubK0j  )��}�(h�h�j  ]�j  K%j  K0ubK1j  )��}�(h�h�j  ]�j  K%j  K1ubK2j  )��}�(h�h�j  ]�j  K%j  K2ubK3j  )��}�(h�h�j  ]�j  K%j  K3ubK4j  )��}�(h�h�j  ]�j  K%j  K4ubK5j  )��}�(h�h�j  ]�j  K%j  K5ubK6j  )��}�(h�h�j  ]�j  K%j  K6ubK7j  )��}�(h�h�j  ]�j  K%j  K7ubK8j  )��}�(h�h�j  ]�j  K%j  K8ubK9j  )��}�(h�h�j  ]�j  K%j  K9ubK:j  )��}�(h�h�j  ]�j  K%j  K:ubK;j  )��}�(h�h�j  ]�j  K%j  K;ubK<j  )��}�(h�h�j  ]�j  K%j  K<ubK=j  )��}�(h�h�j  ]�j  K%j  K=ubK>j  )��}�(h�h�j  ]�j  K%j  K>ubK?j  )��}�(h�h�j  ]�j  K%j  K?ubK@j  )��}�(h�h�j  ]�j  K%j  K@ubKAj  )��}�(h�h�j  ]�j  K%j  KAubKBj  )��}�(h�h�j  ]�j  K%j  KBubKCj  )��}�(h�h�j  ]�j  K%j  KCubKDj  )��}�(h�h�j  ]�j  K%j  KDubKEj  )��}�(h�h�j  ]�j  K%j  KEubKFj  )��}�(h�h�j  ]�j  K%j  KFubKGj  )��}�(h�h�j  ]�j  K%j  KGubKHj  )��}�(h�h�j  ]�j  K%j  KHubKIj  )��}�(h�h�j  ]�j  K%j  KIubKJj  )��}�(h�h�j  ]�j  K%j  KJubKKj  )��}�(h�h�j  ]�j  K%j  KKubKLj  )��}�(h�h�j  ]�j  K%j  KLubKMj  )��}�(h�h�j  ]�j  K%j  KMubKNj  )��}�(h�h�j  ]�j  K%j  KNubKOj  )��}�(h�h�j  ]�j  K%j  KOubuK&}�(K j  )��}�(h�h�j  ]�j  K&j  K ubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubK	j  )��}�(h�h�j  ]�j  K&j  K	ubK
j  )��}�(h�h�j  ]�j  K&j  K
ubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�K5aj  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubKj  )��}�(h�h�j  ]�j  K&j  KubK j  )��}�(h�h�j  ]�j  K&j  K ubK!j  )��}�(h�h�j  ]�j  K&j  K!ubK"j  )��}�(h�h�j  ]�j  K&j  K"ubK#j  )��}�(h�h�j  ]�j  K&j  K#ubK$j  )��}�(h�h�j  ]�j  K&j  K$ubK%j  )��}�(h�h�j  ]�j  K&j  K%ubK&j  )��}�(h�h�j  ]�j  K&j  K&ubK'j  )��}�(h�h�j  ]�j  K&j  K'ubK(j  )��}�(h�h�j  ]�j  K&j  K(ubK)j  )��}�(h�h�j  ]�j  K&j  K)ubK*j  )��}�(h�h�j  ]�j  K&j  K*ubK+j  )��}�(h�h�j  ]�j  K&j  K+ubK,j  )��}�(h�h�j  ]�j  K&j  K,ubK-j  )��}�(h�h�j  ]�j  K&j  K-ubK.j  )��}�(h�h�j  ]�j  K&j  K.ubK/j  )��}�(h�h�j  ]�j  K&j  K/ubK0j  )��}�(h�h�j  ]�j  K&j  K0ubK1j  )��}�(h�h�j  ]�j  K&j  K1ubK2j  )��}�(h�h�j  ]�j  K&j  K2ubK3j  )��}�(h�h�j  ]�j  K&j  K3ubK4j  )��}�(h�h�j  ]�j  K&j  K4ubK5j  )��}�(h�h�j  ]�j  K&j  K5ubK6j  )��}�(h�h�j  ]�j  K&j  K6ubK7j  )��}�(h�h�j  ]�j  K&j  K7ubK8j  )��}�(h�h�j  ]�j  K&j  K8ubK9j  )��}�(h�h�j  ]�j  K&j  K9ubK:j  )��}�(h�h�j  ]�j  K&j  K:ubK;j  )��}�(h�h�j  ]�j  K&j  K;ubK<j  )��}�(h�h�j  ]�j  K&j  K<ubK=j  )��}�(h�h�j  ]�j  K&j  K=ubK>j  )��}�(h�h�j  ]�j  K&j  K>ubK?j  )��}�(h�h�j  ]�j  K&j  K?ubK@j  )��}�(h�h�j  ]�j  K&j  K@ubKAj  )��}�(h�h�j  ]�j  K&j  KAubKBj  )��}�(h�h�j  ]�j  K&j  KBubKCj  )��}�(h�h�j  ]�j  K&j  KCubKDj  )��}�(h�h�j  ]�j  K&j  KDubKEj  )��}�(h�h�j  ]�j  K&j  KEubKFj  )��}�(h�h�j  ]�j  K&j  KFubKGj  )��}�(h�h�j  ]�j  K&j  KGubKHj  )��}�(h�h�j  ]�j  K&j  KHubKIj  )��}�(h�h�j  ]�j  K&j  KIubKJj  )��}�(h�h�j  ]�j  K&j  KJubKKj  )��}�(h�h�j  ]�j  K&j  KKubKLj  )��}�(h�h�j  ]�j  K&j  KLubKMj  )��}�(h�h�j  ]�j  K&j  KMubKNj  )��}�(h�h�j  ]�j  K&j  KNubKOj  )��}�(h�h�j  ]�j  K&j  KOubuK'}�(K j  )��}�(h�h�j  ]�j  K'j  K ubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubK	j  )��}�(h�h�j  ]�j  K'j  K	ubK
j  )��}�(h�h�j  ]�j  K'j  K
ubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubKj  )��}�(h�h�j  ]�j  K'j  KubK j  )��}�(h�h�j  ]�j  K'j  K ubK!j  )��}�(h�h�j  ]�j  K'j  K!ubK"j  )��}�(h�h�j  ]�j  K'j  K"ubK#j  )��}�(h�h�j  ]�j  K'j  K#ubK$j  )��}�(h�h�j  ]�j  K'j  K$ubK%j  )��}�(h�h�j  ]�j  K'j  K%ubK&j  )��}�(h�h�j  ]�j  K'j  K&ubK'j  )��}�(h�h�j  ]�j  K'j  K'ubK(j  )��}�(h�h�j  ]�j  K'j  K(ubK)j  )��}�(h�h�j  ]�j  K'j  K)ubK*j  )��}�(h�h�j  ]�j  K'j  K*ubK+j  )��}�(h�h�j  ]�j  K'j  K+ubK,j  )��}�(h�h�j  ]�j  K'j  K,ubK-j  )��}�(h�h�j  ]�j  K'j  K-ubK.j  )��}�(h�h�j  ]�j  K'j  K.ubK/j  )��}�(h�h�j  ]�j  K'j  K/ubK0j  )��}�(h�h�j  ]�j  K'j  K0ubK1j  )��}�(h�h�j  ]�j  K'j  K1ubK2j  )��}�(h�h�j  ]�j  K'j  K2ubK3j  )��}�(h�h�j  ]�j  K'j  K3ubK4j  )��}�(h�h�j  ]�j  K'j  K4ubK5j  )��}�(h�h�j  ]�j  K'j  K5ubK6j  )��}�(h�h�j  ]�j  K'j  K6ubK7j  )��}�(h�h�j  ]�j  K'j  K7ubK8j  )��}�(h�h�j  ]�j  K'j  K8ubK9j  )��}�(h�h�j  ]�j  K'j  K9ubK:j  )��}�(h�h�j  ]�j  K'j  K:ubK;j  )��}�(h�h�j  ]�j  K'j  K;ubK<j  )��}�(h�h�j  ]�j  K'j  K<ubK=j  )��}�(h�h�j  ]�j  K'j  K=ubK>j  )��}�(h�h�j  ]�j  K'j  K>ubK?j  )��}�(h�h�j  ]�j  K'j  K?ubK@j  )��}�(h�h�j  ]�j  K'j  K@ubKAj  )��}�(h�h�j  ]�j  K'j  KAubKBj  )��}�(h�h�j  ]�j  K'j  KBubKCj  )��}�(h�h�j  ]�j  K'j  KCubKDj  )��}�(h�h�j  ]�j  K'j  KDubKEj  )��}�(h�h�j  ]�j  K'j  KEubKFj  )��}�(h�h�j  ]�j  K'j  KFubKGj  )��}�(h�h�j  ]�j  K'j  KGubKHj  )��}�(h�h�j  ]�j  K'j  KHubKIj  )��}�(h�h�j  ]�j  K'j  KIubKJj  )��}�(h�h�j  ]�j  K'j  KJubKKj  )��}�(h�h�j  ]�j  K'j  KKubKLj  )��}�(h�h�j  ]�j  K'j  KLubKMj  )��}�(h�h�j  ]�j  K'j  KMubKNj  )��}�(h�h�j  ]�j  K'j  KNubKOj  )��}�(h�h�j  ]�j  K'j  KOubuK(}�(K j  )��}�(h�h�j  ]�j  K(j  K ubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubK	j  )��}�(h�h�j  ]�j  K(j  K	ubK
j  )��}�(h�h�j  ]�j  K(j  K
ubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubKj  )��}�(h�h�j  ]�j  K(j  KubK j  )��}�(h�h�j  ]�j  K(j  K ubK!j  )��}�(h�h�j  ]�j  K(j  K!ubK"j  )��}�(h�h�j  ]�j  K(j  K"ubK#j  )��}�(h�h�j  ]�j  K(j  K#ubK$j  )��}�(h�h�j  ]�j  K(j  K$ubK%j  )��}�(h�h�j  ]�j  K(j  K%ubK&j  )��}�(h�h�j  ]�j  K(j  K&ubK'j  )��}�(h�h�j  ]�j  K(j  K'ubK(j  )��}�(h�h�j  ]�j  K(j  K(ubK)j  )��}�(h�h�j  ]�j  K(j  K)ubK*j  )��}�(h�h�j  ]�j  K(j  K*ubK+j  )��}�(h�h�j  ]�j  K(j  K+ubK,j  )��}�(h�h�j  ]�j  K(j  K,ubK-j  )��}�(h�h�j  ]�j  K(j  K-ubK.j  )��}�(h�h�j  ]�j  K(j  K.ubK/j  )��}�(h�h�j  ]�j  K(j  K/ubK0j  )��}�(h�h�j  ]�j  K(j  K0ubK1j  )��}�(h�h�j  ]�j  K(j  K1ubK2j  )��}�(h�h�j  ]�j  K(j  K2ubK3j  )��}�(h�h�j  ]�j  K(j  K3ubK4j  )��}�(h�h�j  ]�j  K(j  K4ubK5j  )��}�(h�h�j  ]�j  K(j  K5ubK6j  )��}�(h�h�j  ]�j  K(j  K6ubK7j  )��}�(h�h�j  ]�j  K(j  K7ubK8j  )��}�(h�h�j  ]�j  K(j  K8ubK9j  )��}�(h�h�j  ]�j  K(j  K9ubK:j  )��}�(h�h�j  ]�j  K(j  K:ubK;j  )��}�(h�h�j  ]�j  K(j  K;ubK<j  )��}�(h�h�j  ]�j  K(j  K<ubK=j  )��}�(h�h�j  ]�j  K(j  K=ubK>j  )��}�(h�h�j  ]�j  K(j  K>ubK?j  )��}�(h�h�j  ]�j  K(j  K?ubK@j  )��}�(h�h�j  ]�j  K(j  K@ubKAj  )��}�(h�h�j  ]�j  K(j  KAubKBj  )��}�(h�h�j  ]�j  K(j  KBubKCj  )��}�(h�h�j  ]�j  K(j  KCubKDj  )��}�(h�h�j  ]�j  K(j  KDubKEj  )��}�(h�h�j  ]�j  K(j  KEubKFj  )��}�(h�h�j  ]�j  K(j  KFubKGj  )��}�(h�h�j  ]�j  K(j  KGubKHj  )��}�(h�h�j  ]�j  K(j  KHubKIj  )��}�(h�h�j  ]�j  K(j  KIubKJj  )��}�(h�h�j  ]�j  K(j  KJubKKj  )��}�(h�h�j  ]�j  K(j  KKubKLj  )��}�(h�h�j  ]�j  K(j  KLubKMj  )��}�(h�h�j  ]�j  K(j  KMubKNj  )��}�(h�h�j  ]�j  K(j  KNubKOj  )��}�(h�h�j  ]�j  K(j  KOubuK)}�(K j  )��}�(h�h�j  ]�j  K)j  K ubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubK	j  )��}�(h�h�j  ]�j  K)j  K	ubK
j  )��}�(h�h�j  ]�j  K)j  K
ubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubKj  )��}�(h�h�j  ]�j  K)j  KubK j  )��}�(h�h�j  ]�j  K)j  K ubK!j  )��}�(h�h�j  ]�j  K)j  K!ubK"j  )��}�(h�h�j  ]�j  K)j  K"ubK#j  )��}�(h�h�j  ]�j  K)j  K#ubK$j  )��}�(h�h�j  ]�j  K)j  K$ubK%j  )��}�(h�h�j  ]�j  K)j  K%ubK&j  )��}�(h�h�j  ]�j  K)j  K&ubK'j  )��}�(h�h�j  ]�j  K)j  K'ubK(j  )��}�(h�h�j  ]�j  K)j  K(ubK)j  )��}�(h�h�j  ]�j  K)j  K)ubK*j  )��}�(h�h�j  ]�j  K)j  K*ubK+j  )��}�(h�h�j  ]�j  K)j  K+ubK,j  )��}�(h�h�j  ]�j  K)j  K,ubK-j  )��}�(h�h�j  ]�j  K)j  K-ubK.j  )��}�(h�h�j  ]�j  K)j  K.ubK/j  )��}�(h�h�j  ]�j  K)j  K/ubK0j  )��}�(h�h�j  ]�j  K)j  K0ubK1j  )��}�(h�h�j  ]�j  K)j  K1ubK2j  )��}�(h�h�j  ]�j  K)j  K2ubK3j  )��}�(h�h�j  ]�j  K)j  K3ubK4j  )��}�(h�h�j  ]�j  K)j  K4ubK5j  )��}�(h�h�j  ]�j  K)j  K5ubK6j  )��}�(h�h�j  ]�j  K)j  K6ubK7j  )��}�(h�h�j  ]�j  K)j  K7ubK8j  )��}�(h�h�j  ]�j  K)j  K8ubK9j  )��}�(h�h�j  ]�j  K)j  K9ubK:j  )��}�(h�h�j  ]�j  K)j  K:ubK;j  )��}�(h�h�j  ]�j  K)j  K;ubK<j  )��}�(h�h�j  ]�j  K)j  K<ubK=j  )��}�(h�h�j  ]�j  K)j  K=ubK>j  )��}�(h�h�j  ]�j  K)j  K>ubK?j  )��}�(h�h�j  ]�j  K)j  K?ubK@j  )��}�(h�h�j  ]�j  K)j  K@ubKAj  )��}�(h�h�j  ]�j  K)j  KAubKBj  )��}�(h�h�j  ]�j  K)j  KBubKCj  )��}�(h�h�j  ]�j  K)j  KCubKDj  )��}�(h�h�j  ]�j  K)j  KDubKEj  )��}�(h�h�j  ]�j  K)j  KEubKFj  )��}�(h�h�j  ]�j  K)j  KFubKGj  )��}�(h�h�j  ]�j  K)j  KGubKHj  )��}�(h�h�j  ]�j  K)j  KHubKIj  )��}�(h�h�j  ]�j  K)j  KIubKJj  )��}�(h�h�j  ]�j  K)j  KJubKKj  )��}�(h�h�j  ]�j  K)j  KKubKLj  )��}�(h�h�j  ]�j  K)j  KLubKMj  )��}�(h�h�j  ]�j  K)j  KMubKNj  )��}�(h�h�j  ]�j  K)j  KNubKOj  )��}�(h�h�j  ]�j  K)j  KOubuK*}�(K j  )��}�(h�h�j  ]�j  K*j  K ubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubK	j  )��}�(h�h�j  ]�j  K*j  K	ubK
j  )��}�(h�h�j  ]�j  K*j  K
ubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubKj  )��}�(h�h�j  ]�j  K*j  KubK j  )��}�(h�h�j  ]�j  K*j  K ubK!j  )��}�(h�h�j  ]�j  K*j  K!ubK"j  )��}�(h�h�j  ]�j  K*j  K"ubK#j  )��}�(h�h�j  ]�j  K*j  K#ubK$j  )��}�(h�h�j  ]�j  K*j  K$ubK%j  )��}�(h�h�j  ]�j  K*j  K%ubK&j  )��}�(h�h�j  ]�j  K*j  K&ubK'j  )��}�(h�h�j  ]�j  K*j  K'ubK(j  )��}�(h�h�j  ]�j  K*j  K(ubK)j  )��}�(h�h�j  ]�j  K*j  K)ubK*j  )��}�(h�h�j  ]�j  K*j  K*ubK+j  )��}�(h�h�j  ]�j  K*j  K+ubK,j  )��}�(h�h�j  ]�j  K*j  K,ubK-j  )��}�(h�h�j  ]�j  K*j  K-ubK.j  )��}�(h�h�j  ]�j  K*j  K.ubK/j  )��}�(h�h�j  ]�j  K*j  K/ubK0j  )��}�(h�h�j  ]�j  K*j  K0ubK1j  )��}�(h�h�j  ]�j  K*j  K1ubK2j  )��}�(h�h�j  ]�j  K*j  K2ubK3j  )��}�(h�h�j  ]�j  K*j  K3ubK4j  )��}�(h�h�j  ]�j  K*j  K4ubK5j  )��}�(h�h�j  ]�j  K*j  K5ubK6j  )��}�(h�h�j  ]�j  K*j  K6ubK7j  )��}�(h�h�j  ]�j  K*j  K7ubK8j  )��}�(h�h�j  ]�j  K*j  K8ubK9j  )��}�(h�h�j  ]�j  K*j  K9ubK:j  )��}�(h�h�j  ]�j  K*j  K:ubK;j  )��}�(h�h�j  ]�j  K*j  K;ubK<j  )��}�(h�h�j  ]�j  K*j  K<ubK=j  )��}�(h�h�j  ]�j  K*j  K=ubK>j  )��}�(h�h�j  ]�j  K*j  K>ubK?j  )��}�(h�h�j  ]�j  K*j  K?ubK@j  )��}�(h�h�j  ]�j  K*j  K@ubKAj  )��}�(h�h�j  ]�j  K*j  KAubKBj  )��}�(h�h�j  ]�j  K*j  KBubKCj  )��}�(h�h�j  ]�j  K*j  KCubKDj  )��}�(h�h�j  ]�j  K*j  KDubKEj  )��}�(h�h�j  ]�j  K*j  KEubKFj  )��}�(h�h�j  ]�j  K*j  KFubKGj  )��}�(h�h�j  ]�j  K*j  KGubKHj  )��}�(h�h�j  ]�j  K*j  KHubKIj  )��}�(h�h�j  ]�j  K*j  KIubKJj  )��}�(h�h�j  ]�j  K*j  KJubKKj  )��}�(h�h�j  ]�j  K*j  KKubKLj  )��}�(h�h�j  ]�j  K*j  KLubKMj  )��}�(h�h�j  ]�j  K*j  KMubKNj  )��}�(h�h�j  ]�j  K*j  KNubKOj  )��}�(h�h�j  ]�j  K*j  KOubuK+}�(K j  )��}�(h�h�j  ]�j  K+j  K ubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubK	j  )��}�(h�h�j  ]�j  K+j  K	ubK
j  )��}�(h�h�j  ]�j  K+j  K
ubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubKj  )��}�(h�h�j  ]�j  K+j  KubK j  )��}�(h�h�j  ]�j  K+j  K ubK!j  )��}�(h�h�j  ]�j  K+j  K!ubK"j  )��}�(h�h�j  ]�j  K+j  K"ubK#j  )��}�(h�h�j  ]�j  K+j  K#ubK$j  )��}�(h�h�j  ]�j  K+j  K$ubK%j  )��}�(h�h�j  ]�j  K+j  K%ubK&j  )��}�(h�h�j  ]�j  K+j  K&ubK'j  )��}�(h�h�j  ]�j  K+j  K'ubK(j  )��}�(h�h�j  ]�j  K+j  K(ubK)j  )��}�(h�h�j  ]�j  K+j  K)ubK*j  )��}�(h�h�j  ]�j  K+j  K*ubK+j  )��}�(h�h�j  ]�j  K+j  K+ubK,j  )��}�(h�h�j  ]�j  K+j  K,ubK-j  )��}�(h�h�j  ]�j  K+j  K-ubK.j  )��}�(h�h�j  ]�j  K+j  K.ubK/j  )��}�(h�h�j  ]�j  K+j  K/ubK0j  )��}�(h�h�j  ]�j  K+j  K0ubK1j  )��}�(h�h�j  ]�j  K+j  K1ubK2j  )��}�(h�h�j  ]�j  K+j  K2ubK3j  )��}�(h�h�j  ]�j  K+j  K3ubK4j  )��}�(h�h�j  ]�j  K+j  K4ubK5j  )��}�(h�h�j  ]�j  K+j  K5ubK6j  )��}�(h�h�j  ]�j  K+j  K6ubK7j  )��}�(h�h�j  ]�j  K+j  K7ubK8j  )��}�(h�h�j  ]�j  K+j  K8ubK9j  )��}�(h�h�j  ]�j  K+j  K9ubK:j  )��}�(h�h�j  ]�j  K+j  K:ubK;j  )��}�(h�h�j  ]�j  K+j  K;ubK<j  )��}�(h�h�j  ]�j  K+j  K<ubK=j  )��}�(h�h�j  ]�j  K+j  K=ubK>j  )��}�(h�h�j  ]�j  K+j  K>ubK?j  )��}�(h�h�j  ]�j  K+j  K?ubK@j  )��}�(h�h�j  ]�j  K+j  K@ubKAj  )��}�(h�h�j  ]�j  K+j  KAubKBj  )��}�(h�h�j  ]�j  K+j  KBubKCj  )��}�(h�h�j  ]�j  K+j  KCubKDj  )��}�(h�h�j  ]�j  K+j  KDubKEj  )��}�(h�h�j  ]�j  K+j  KEubKFj  )��}�(h�h�j  ]�j  K+j  KFubKGj  )��}�(h�h�j  ]�j  K+j  KGubKHj  )��}�(h�h�j  ]�j  K+j  KHubKIj  )��}�(h�h�j  ]�j  K+j  KIubKJj  )��}�(h�h�j  ]�j  K+j  KJubKKj  )��}�(h�h�j  ]�j  K+j  KKubKLj  )��}�(h�h�j  ]�j  K+j  KLubKMj  )��}�(h�h�j  ]�j  K+j  KMubKNj  )��}�(h�h�j  ]�j  K+j  KNubKOj  )��}�(h�h�j  ]�j  K+j  KOubuK,}�(K j  )��}�(h�h�j  ]�j  K,j  K ubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubK	j  )��}�(h�h�j  ]�j  K,j  K	ubK
j  )��}�(h�h�j  ]�j  K,j  K
ubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubKj  )��}�(h�h�j  ]�j  K,j  KubK j  )��}�(h�h�j  ]�j  K,j  K ubK!j  )��}�(h�h�j  ]�j  K,j  K!ubK"j  )��}�(h�h�j  ]�j  K,j  K"ubK#j  )��}�(h�h�j  ]�j  K,j  K#ubK$j  )��}�(h�h�j  ]�j  K,j  K$ubK%j  )��}�(h�h�j  ]�j  K,j  K%ubK&j  )��}�(h�h�j  ]�j  K,j  K&ubK'j  )��}�(h�h�j  ]�j  K,j  K'ubK(j  )��}�(h�h�j  ]�j  K,j  K(ubK)j  )��}�(h�h�j  ]�j  K,j  K)ubK*j  )��}�(h�h�j  ]�j  K,j  K*ubK+j  )��}�(h�h�j  ]�j  K,j  K+ubK,j  )��}�(h�h�j  ]�j  K,j  K,ubK-j  )��}�(h�h�j  ]�j  K,j  K-ubK.j  )��}�(h�h�j  ]�j  K,j  K.ubK/j  )��}�(h�h�j  ]�j  K,j  K/ubK0j  )��}�(h�h�j  ]�j  K,j  K0ubK1j  )��}�(h�h�j  ]�j  K,j  K1ubK2j  )��}�(h�h�j  ]�j  K,j  K2ubK3j  )��}�(h�h�j  ]�j  K,j  K3ubK4j  )��}�(h�h�j  ]�j  K,j  K4ubK5j  )��}�(h�h�j  ]�j  K,j  K5ubK6j  )��}�(h�h�j  ]�j  K,j  K6ubK7j  )��}�(h�h�j  ]�j  K,j  K7ubK8j  )��}�(h�h�j  ]�j  K,j  K8ubK9j  )��}�(h�h�j  ]�j  K,j  K9ubK:j  )��}�(h�h�j  ]�j  K,j  K:ubK;j  )��}�(h�h�j  ]�j  K,j  K;ubK<j  )��}�(h�h�j  ]�j  K,j  K<ubK=j  )��}�(h�h�j  ]�j  K,j  K=ubK>j  )��}�(h�h�j  ]�j  K,j  K>ubK?j  )��}�(h�h�j  ]�j  K,j  K?ubK@j  )��}�(h�h�j  ]�j  K,j  K@ubKAj  )��}�(h�h�j  ]�j  K,j  KAubKBj  )��}�(h�h�j  ]�j  K,j  KBubKCj  )��}�(h�h�j  ]�j  K,j  KCubKDj  )��}�(h�h�j  ]�j  K,j  KDubKEj  )��}�(h�h�j  ]�j  K,j  KEubKFj  )��}�(h�h�j  ]�j  K,j  KFubKGj  )��}�(h�h�j  ]�j  K,j  KGubKHj  )��}�(h�h�j  ]�j  K,j  KHubKIj  )��}�(h�h�j  ]�j  K,j  KIubKJj  )��}�(h�h�j  ]�j  K,j  KJubKKj  )��}�(h�h�j  ]�j  K,j  KKubKLj  )��}�(h�h�j  ]�j  K,j  KLubKMj  )��}�(h�h�j  ]�j  K,j  KMubKNj  )��}�(h�h�j  ]�j  K,j  KNubKOj  )��}�(h�h�j  ]�j  K,j  KOubuK-}�(K j  )��}�(h�h�j  ]�j  K-j  K ubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubK	j  )��}�(h�h�j  ]�j  K-j  K	ubK
j  )��}�(h�h�j  ]�j  K-j  K
ubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubKj  )��}�(h�h�j  ]�j  K-j  KubK j  )��}�(h�h�j  ]�j  K-j  K ubK!j  )��}�(h�h�j  ]�j  K-j  K!ubK"j  )��}�(h�h�j  ]�j  K-j  K"ubK#j  )��}�(h�h�j  ]�j  K-j  K#ubK$j  )��}�(h�h�j  ]�j  K-j  K$ubK%j  )��}�(h�h�j  ]�j  K-j  K%ubK&j  )��}�(h�h�j  ]�j  K-j  K&ubK'j  )��}�(h�h�j  ]�j  K-j  K'ubK(j  )��}�(h�h�j  ]�j  K-j  K(ubK)j  )��}�(h�h�j  ]�j  K-j  K)ubK*j  )��}�(h�h�j  ]�j  K-j  K*ubK+j  )��}�(h�h�j  ]�j  K-j  K+ubK,j  )��}�(h�h�j  ]�j  K-j  K,ubK-j  )��}�(h�h�j  ]�j  K-j  K-ubK.j  )��}�(h�h�j  ]�j  K-j  K.ubK/j  )��}�(h�h�j  ]�j  K-j  K/ubK0j  )��}�(h�h�j  ]�j  K-j  K0ubK1j  )��}�(h�h�j  ]�j  K-j  K1ubK2j  )��}�(h�h�j  ]�j  K-j  K2ubK3j  )��}�(h�h�j  ]�j  K-j  K3ubK4j  )��}�(h�h�j  ]�j  K-j  K4ubK5j  )��}�(h�h�j  ]�j  K-j  K5ubK6j  )��}�(h�h�j  ]�j  K-j  K6ubK7j  )��}�(h�h�j  ]�j  K-j  K7ubK8j  )��}�(h�h�j  ]�j  K-j  K8ubK9j  )��}�(h�h�j  ]�j  K-j  K9ubK:j  )��}�(h�h�j  ]�j  K-j  K:ubK;j  )��}�(h�h�j  ]�j  K-j  K;ubK<j  )��}�(h�h�j  ]�j  K-j  K<ubK=j  )��}�(h�h�j  ]�j  K-j  K=ubK>j  )��}�(h�h�j  ]�j  K-j  K>ubK?j  )��}�(h�h�j  ]�j  K-j  K?ubK@j  )��}�(h�h�j  ]�j  K-j  K@ubKAj  )��}�(h�h�j  ]�j  K-j  KAubKBj  )��}�(h�h�j  ]�j  K-j  KBubKCj  )��}�(h�h�j  ]�j  K-j  KCubKDj  )��}�(h�h�j  ]�j  K-j  KDubKEj  )��}�(h�h�j  ]�j  K-j  KEubKFj  )��}�(h�h�j  ]�j  K-j  KFubKGj  )��}�(h�h�j  ]�j  K-j  KGubKHj  )��}�(h�h�j  ]�j  K-j  KHubKIj  )��}�(h�h�j  ]�j  K-j  KIubKJj  )��}�(h�h�j  ]�j  K-j  KJubKKj  )��}�(h�h�j  ]�j  K-j  KKubKLj  )��}�(h�h�j  ]�j  K-j  KLubKMj  )��}�(h�h�j  ]�j  K-j  KMubKNj  )��}�(h�h�j  ]�j  K-j  KNubKOj  )��}�(h�h�j  ]�j  K-j  KOubuK.}�(K j  )��}�(h�h�j  ]�j  K.j  K ubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubK	j  )��}�(h�h�j  ]�j  K.j  K	ubK
j  )��}�(h�h�j  ]�j  K.j  K
ubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubKj  )��}�(h�h�j  ]�j  K.j  KubK j  )��}�(h�h�j  ]�j  K.j  K ubK!j  )��}�(h�h�j  ]�j  K.j  K!ubK"j  )��}�(h�h�j  ]�j  K.j  K"ubK#j  )��}�(h�h�j  ]�j  K.j  K#ubK$j  )��}�(h�h�j  ]�j  K.j  K$ubK%j  )��}�(h�h�j  ]�j  K.j  K%ubK&j  )��}�(h�h�j  ]�j  K.j  K&ubK'j  )��}�(h�h�j  ]�j  K.j  K'ubK(j  )��}�(h�h�j  ]�j  K.j  K(ubK)j  )��}�(h�h�j  ]�j  K.j  K)ubK*j  )��}�(h�h�j  ]�j  K.j  K*ubK+j  )��}�(h�h�j  ]�j  K.j  K+ubK,j  )��}�(h�h�j  ]�j  K.j  K,ubK-j  )��}�(h�h�j  ]�j  K.j  K-ubK.j  )��}�(h�h�j  ]�j  K.j  K.ubK/j  )��}�(h�h�j  ]�j  K.j  K/ubK0j  )��}�(h�h�j  ]�j  K.j  K0ubK1j  )��}�(h�h�j  ]�j  K.j  K1ubK2j  )��}�(h�h�j  ]�j  K.j  K2ubK3j  )��}�(h�h�j  ]�j  K.j  K3ubK4j  )��}�(h�h�j  ]�j  K.j  K4ubK5j  )��}�(h�h�j  ]�j  K.j  K5ubK6j  )��}�(h�h�j  ]�j  K.j  K6ubK7j  )��}�(h�h�j  ]�j  K.j  K7ubK8j  )��}�(h�h�j  ]�j  K.j  K8ubK9j  )��}�(h�h�j  ]�j  K.j  K9ubK:j  )��}�(h�h�j  ]�j  K.j  K:ubK;j  )��}�(h�h�j  ]�j  K.j  K;ubK<j  )��}�(h�h�j  ]�j  K.j  K<ubK=j  )��}�(h�h�j  ]�j  K.j  K=ubK>j  )��}�(h�h�j  ]�j  K.j  K>ubK?j  )��}�(h�h�j  ]�j  K.j  K?ubK@j  )��}�(h�h�j  ]�j  K.j  K@ubKAj  )��}�(h�h�j  ]�j  K.j  KAubKBj  )��}�(h�h�j  ]�j  K.j  KBubKCj  )��}�(h�h�j  ]�j  K.j  KCubKDj  )��}�(h�h�j  ]�j  K.j  KDubKEj  )��}�(h�h�j  ]�j  K.j  KEubKFj  )��}�(h�h�j  ]�j  K.j  KFubKGj  )��}�(h�h�j  ]�j  K.j  KGubKHj  )��}�(h�h�j  ]�j  K.j  KHubKIj  )��}�(h�h�j  ]�j  K.j  KIubKJj  )��}�(h�h�j  ]�j  K.j  KJubKKj  )��}�(h�h�j  ]�j  K.j  KKubKLj  )��}�(h�h�j  ]�j  K.j  KLubKMj  )��}�(h�h�j  ]�j  K.j  KMubKNj  )��}�(h�h�j  ]�j  K.j  KNubKOj  )��}�(h�h�j  ]�j  K.j  KOubuK/}�(K j  )��}�(h�h�j  ]�j  K/j  K ubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubK	j  )��}�(h�h�j  ]�j  K/j  K	ubK
j  )��}�(h�h�j  ]�j  K/j  K
ubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubKj  )��}�(h�h�j  ]�j  K/j  KubK j  )��}�(h�h�j  ]�j  K/j  K ubK!j  )��}�(h�h�j  ]�j  K/j  K!ubK"j  )��}�(h�h�j  ]�j  K/j  K"ubK#j  )��}�(h�h�j  ]�j  K/j  K#ubK$j  )��}�(h�h�j  ]�j  K/j  K$ubK%j  )��}�(h�h�j  ]�j  K/j  K%ubK&j  )��}�(h�h�j  ]�j  K/j  K&ubK'j  )��}�(h�h�j  ]�j  K/j  K'ubK(j  )��}�(h�h�j  ]�j  K/j  K(ubK)j  )��}�(h�h�j  ]�j  K/j  K)ubK*j  )��}�(h�h�j  ]�j  K/j  K*ubK+j  )��}�(h�h�j  ]�j  K/j  K+ubK,j  )��}�(h�h�j  ]�j  K/j  K,ubK-j  )��}�(h�h�j  ]�j  K/j  K-ubK.j  )��}�(h�h�j  ]�j  K/j  K.ubK/j  )��}�(h�h�j  ]�K6aj  K/j  K/ubK0j  )��}�(h�h�j  ]�j  K/j  K0ubK1j  )��}�(h�h�j  ]�j  K/j  K1ubK2j  )��}�(h�h�j  ]�j  K/j  K2ubK3j  )��}�(h�h�j  ]�j  K/j  K3ubK4j  )��}�(h�h�j  ]�j  K/j  K4ubK5j  )��}�(h�h�j  ]�j  K/j  K5ubK6j  )��}�(h�h�j  ]�j  K/j  K6ubK7j  )��}�(h�h�j  ]�j  K/j  K7ubK8j  )��}�(h�h�j  ]�j  K/j  K8ubK9j  )��}�(h�h�j  ]�j  K/j  K9ubK:j  )��}�(h�h�j  ]�j  K/j  K:ubK;j  )��}�(h�h�j  ]�j  K/j  K;ubK<j  )��}�(h�h�j  ]�j  K/j  K<ubK=j  )��}�(h�h�j  ]�j  K/j  K=ubK>j  )��}�(h�h�j  ]�j  K/j  K>ubK?j  )��}�(h�h�j  ]�j  K/j  K?ubK@j  )��}�(h�h�j  ]�j  K/j  K@ubKAj  )��}�(h�h�j  ]�j  K/j  KAubKBj  )��}�(h�h�j  ]�j  K/j  KBubKCj  )��}�(h�h�j  ]�j  K/j  KCubKDj  )��}�(h�h�j  ]�j  K/j  KDubKEj  )��}�(h�h�j  ]�j  K/j  KEubKFj  )��}�(h�h�j  ]�j  K/j  KFubKGj  )��}�(h�h�j  ]�j  K/j  KGubKHj  )��}�(h�h�j  ]�j  K/j  KHubKIj  )��}�(h�h�j  ]�j  K/j  KIubKJj  )��}�(h�h�j  ]�j  K/j  KJubKKj  )��}�(h�h�j  ]�j  K/j  KKubKLj  )��}�(h�h�j  ]�j  K/j  KLubKMj  )��}�(h�h�j  ]�j  K/j  KMubKNj  )��}�(h�h�j  ]�j  K/j  KNubKOj  )��}�(h�h�j  ]�j  K/j  KOubuK0}�(K j  )��}�(h�h�j  ]�j  K0j  K ubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubK	j  )��}�(h�h�j  ]�j  K0j  K	ubK
j  )��}�(h�h�j  ]�j  K0j  K
ubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubKj  )��}�(h�h�j  ]�j  K0j  KubK j  )��}�(h�h�j  ]�j  K0j  K ubK!j  )��}�(h�h�j  ]�j  K0j  K!ubK"j  )��}�(h�h�j  ]�j  K0j  K"ubK#j  )��}�(h�h�j  ]�j  K0j  K#ubK$j  )��}�(h�h�j  ]�j  K0j  K$ubK%j  )��}�(h�h�j  ]�j  K0j  K%ubK&j  )��}�(h�h�j  ]�j  K0j  K&ubK'j  )��}�(h�h�j  ]�j  K0j  K'ubK(j  )��}�(h�h�j  ]�j  K0j  K(ubK)j  )��}�(h�h�j  ]�j  K0j  K)ubK*j  )��}�(h�h�j  ]�K8aj  K0j  K*ubK+j  )��}�(h�h�j  ]�j  K0j  K+ubK,j  )��}�(h�h�j  ]�j  K0j  K,ubK-j  )��}�(h�h�j  ]�j  K0j  K-ubK.j  )��}�(h�h�j  ]�j  K0j  K.ubK/j  )��}�(h�h�j  ]�j  K0j  K/ubK0j  )��}�(h�h�j  ]�j  K0j  K0ubK1j  )��}�(h�h�j  ]�j  K0j  K1ubK2j  )��}�(h�h�j  ]�j  K0j  K2ubK3j  )��}�(h�h�j  ]�j  K0j  K3ubK4j  )��}�(h�h�j  ]�j  K0j  K4ubK5j  )��}�(h�h�j  ]�j  K0j  K5ubK6j  )��}�(h�h�j  ]�j  K0j  K6ubK7j  )��}�(h�h�j  ]�j  K0j  K7ubK8j  )��}�(h�h�j  ]�j  K0j  K8ubK9j  )��}�(h�h�j  ]�j  K0j  K9ubK:j  )��}�(h�h�j  ]�j  K0j  K:ubK;j  )��}�(h�h�j  ]�j  K0j  K;ubK<j  )��}�(h�h�j  ]�j  K0j  K<ubK=j  )��}�(h�h�j  ]�j  K0j  K=ubK>j  )��}�(h�h�j  ]�j  K0j  K>ubK?j  )��}�(h�h�j  ]�j  K0j  K?ubK@j  )��}�(h�h�j  ]�j  K0j  K@ubKAj  )��}�(h�h�j  ]�j  K0j  KAubKBj  )��}�(h�h�j  ]�j  K0j  KBubKCj  )��}�(h�h�j  ]�j  K0j  KCubKDj  )��}�(h�h�j  ]�j  K0j  KDubKEj  )��}�(h�h�j  ]�j  K0j  KEubKFj  )��}�(h�h�j  ]�j  K0j  KFubKGj  )��}�(h�h�j  ]�j  K0j  KGubKHj  )��}�(h�h�j  ]�j  K0j  KHubKIj  )��}�(h�h�j  ]�j  K0j  KIubKJj  )��}�(h�h�j  ]�j  K0j  KJubKKj  )��}�(h�h�j  ]�j  K0j  KKubKLj  )��}�(h�h�j  ]�j  K0j  KLubKMj  )��}�(h�h�j  ]�j  K0j  KMubKNj  )��}�(h�h�j  ]�j  K0j  KNubKOj  )��}�(h�h�j  ]�j  K0j  KOubuK1}�(K j  )��}�(h�h�j  ]�j  K1j  K ubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubK	j  )��}�(h�h�j  ]�j  K1j  K	ubK
j  )��}�(h�h�j  ]�j  K1j  K
ubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubKj  )��}�(h�h�j  ]�j  K1j  KubK j  )��}�(h�h�j  ]�j  K1j  K ubK!j  )��}�(h�h�j  ]�j  K1j  K!ubK"j  )��}�(h�h�j  ]�j  K1j  K"ubK#j  )��}�(h�h�j  ]�j  K1j  K#ubK$j  )��}�(h�h�j  ]�j  K1j  K$ubK%j  )��}�(h�h�j  ]�j  K1j  K%ubK&j  )��}�(h�h�j  ]�j  K1j  K&ubK'j  )��}�(h�h�j  ]�j  K1j  K'ubK(j  )��}�(h�h�j  ]�j  K1j  K(ubK)j  )��}�(h�h�j  ]�j  K1j  K)ubK*j  )��}�(h�h�j  ]�j  K1j  K*ubK+j  )��}�(h�h�j  ]�j  K1j  K+ubK,j  )��}�(h�h�j  ]�j  K1j  K,ubK-j  )��}�(h�h�j  ]�j  K1j  K-ubK.j  )��}�(h�h�j  ]�j  K1j  K.ubK/j  )��}�(h�h�j  ]�j  K1j  K/ubK0j  )��}�(h�h�j  ]�j  K1j  K0ubK1j  )��}�(h�h�j  ]�j  K1j  K1ubK2j  )��}�(h�h�j  ]�j  K1j  K2ubK3j  )��}�(h�h�j  ]�j  K1j  K3ubK4j  )��}�(h�h�j  ]�j  K1j  K4ubK5j  )��}�(h�h�j  ]�j  K1j  K5ubK6j  )��}�(h�h�j  ]�j  K1j  K6ubK7j  )��}�(h�h�j  ]�j  K1j  K7ubK8j  )��}�(h�h�j  ]�j  K1j  K8ubK9j  )��}�(h�h�j  ]�j  K1j  K9ubK:j  )��}�(h�h�j  ]�j  K1j  K:ubK;j  )��}�(h�h�j  ]�j  K1j  K;ubK<j  )��}�(h�h�j  ]�j  K1j  K<ubK=j  )��}�(h�h�j  ]�j  K1j  K=ubK>j  )��}�(h�h�j  ]�j  K1j  K>ubK?j  )��}�(h�h�j  ]�j  K1j  K?ubK@j  )��}�(h�h�j  ]�j  K1j  K@ubKAj  )��}�(h�h�j  ]�j  K1j  KAubKBj  )��}�(h�h�j  ]�j  K1j  KBubKCj  )��}�(h�h�j  ]�j  K1j  KCubKDj  )��}�(h�h�j  ]�j  K1j  KDubKEj  )��}�(h�h�j  ]�j  K1j  KEubKFj  )��}�(h�h�j  ]�j  K1j  KFubKGj  )��}�(h�h�j  ]�j  K1j  KGubKHj  )��}�(h�h�j  ]�j  K1j  KHubKIj  )��}�(h�h�j  ]�j  K1j  KIubKJj  )��}�(h�h�j  ]�j  K1j  KJubKKj  )��}�(h�h�j  ]�j  K1j  KKubKLj  )��}�(h�h�j  ]�j  K1j  KLubKMj  )��}�(h�h�j  ]�j  K1j  KMubKNj  )��}�(h�h�j  ]�j  K1j  KNubKOj  )��}�(h�h�j  ]�j  K1j  KOubuK2}�(K j  )��}�(h�h�j  ]�j  K2j  K ubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubK	j  )��}�(h�h�j  ]�j  K2j  K	ubK
j  )��}�(h�h�j  ]�j  K2j  K
ubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubKj  )��}�(h�h�j  ]�j  K2j  KubK j  )��}�(h�h�j  ]�j  K2j  K ubK!j  )��}�(h�h�j  ]�j  K2j  K!ubK"j  )��}�(h�h�j  ]�j  K2j  K"ubK#j  )��}�(h�h�j  ]�j  K2j  K#ubK$j  )��}�(h�h�j  ]�j  K2j  K$ubK%j  )��}�(h�h�j  ]�j  K2j  K%ubK&j  )��}�(h�h�j  ]�j  K2j  K&ubK'j  )��}�(h�h�j  ]�j  K2j  K'ubK(j  )��}�(h�h�j  ]�j  K2j  K(ubK)j  )��}�(h�h�j  ]�j  K2j  K)ubK*j  )��}�(h�h�j  ]�j  K2j  K*ubK+j  )��}�(h�h�j  ]�j  K2j  K+ubK,j  )��}�(h�h�j  ]�j  K2j  K,ubK-j  )��}�(h�h�j  ]�j  K2j  K-ubK.j  )��}�(h�h�j  ]�j  K2j  K.ubK/j  )��}�(h�h�j  ]�j  K2j  K/ubK0j  )��}�(h�h�j  ]�j  K2j  K0ubK1j  )��}�(h�h�j  ]�j  K2j  K1ubK2j  )��}�(h�h�j  ]�j  K2j  K2ubK3j  )��}�(h�h�j  ]�j  K2j  K3ubK4j  )��}�(h�h�j  ]�j  K2j  K4ubK5j  )��}�(h�h�j  ]�j  K2j  K5ubK6j  )��}�(h�h�j  ]�j  K2j  K6ubK7j  )��}�(h�h�j  ]�j  K2j  K7ubK8j  )��}�(h�h�j  ]�j  K2j  K8ubK9j  )��}�(h�h�j  ]�j  K2j  K9ubK:j  )��}�(h�h�j  ]�j  K2j  K:ubK;j  )��}�(h�h�j  ]�j  K2j  K;ubK<j  )��}�(h�h�j  ]�j  K2j  K<ubK=j  )��}�(h�h�j  ]�j  K2j  K=ubK>j  )��}�(h�h�j  ]�j  K2j  K>ubK?j  )��}�(h�h�j  ]�j  K2j  K?ubK@j  )��}�(h�h�j  ]�j  K2j  K@ubKAj  )��}�(h�h�j  ]�j  K2j  KAubKBj  )��}�(h�h�j  ]�j  K2j  KBubKCj  )��}�(h�h�j  ]�j  K2j  KCubKDj  )��}�(h�h�j  ]�j  K2j  KDubKEj  )��}�(h�h�j  ]�j  K2j  KEubKFj  )��}�(h�h�j  ]�j  K2j  KFubKGj  )��}�(h�h�j  ]�j  K2j  KGubKHj  )��}�(h�h�j  ]�j  K2j  KHubKIj  )��}�(h�h�j  ]�j  K2j  KIubKJj  )��}�(h�h�j  ]�j  K2j  KJubKKj  )��}�(h�h�j  ]�j  K2j  KKubKLj  )��}�(h�h�j  ]�j  K2j  KLubKMj  )��}�(h�h�j  ]�j  K2j  KMubKNj  )��}�(h�h�j  ]�j  K2j  KNubKOj  )��}�(h�h�j  ]�j  K2j  KOubuK3}�(K j  )��}�(h�h�j  ]�j  K3j  K ubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubK	j  )��}�(h�h�j  ]�j  K3j  K	ubK
j  )��}�(h�h�j  ]�j  K3j  K
ubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h֕      h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubKj  )��}�(h�h�j  ]�j  K3j  KubK j  )��}�(h�h�j  ]�j  K3j  K ubK!j  )��}�(h�h�j  ]�j  K3j  K!ubK"j  )��}�(h�h�j  ]�j  K3j  K"ubK#j  )��}�(h�h�j  ]�j  K3j  K#ubK$j  )��}�(h�h�j  ]�j  K3j  K$ubK%j  )��}�(h�h�j  ]�j  K3j  K%ubK&j  )��}�(h�h�j  ]�j  K3j  K&ubK'j  )��}�(h�h�j  ]�j  K3j  K'ubK(j  )��}�(h�h�j  ]�j  K3j  K(ubK)j  )��}�(h�h�j  ]�j  K3j  K)ubK*j  )��}�(h�h�j  ]�j  K3j  K*ubK+j  )��}�(h�h�j  ]�j  K3j  K+ubK,j  )��}�(h�h�j  ]�j  K3j  K,ubK-j  )��}�(h�h�j  ]�j  K3j  K-ubK.j  )��}�(h�h�j  ]�j  K3j  K.ubK/j  )��}�(h�h�j  ]�j  K3j  K/ubK0j  )��}�(h�h�j  ]�j  K3j  K0ubK1j  )��}�(h�h�j  ]�j  K3j  K1ubK2j  )��}�(h�h�j  ]�j  K3j  K2ubK3j  )��}�(h�h�j  ]�j  K3j  K3ubK4j  )��}�(h�h�j  ]�j  K3j  K4ubK5j  )��}�(h�h�j  ]�j  K3j  K5ubK6j  )��}�(h�h�j  ]�j  K3j  K6ubK7j  )��}�(h�h�j  ]�j  K3j  K7ubK8j  )��}�(h�h�j  ]�j  K3j  K8ubK9j  )��}�(h�h�j  ]�j  K3j  K9ubK:j  )��}�(h�h�j  ]�j  K3j  K:ubK;j  )��}�(h�h�j  ]�j  K3j  K;ubK<j  )��}�(h�h�j  ]�j  K3j  K<ubK=j  )��}�(h�h�j  ]�j  K3j  K=ubK>j  )��}�(h�h�j  ]�j  K3j  K>ubK?j  )��}�(h�h�j  ]�j  K3j  K?ubK@j  )��}�(h�h�j  ]�j  K3j  K@ubKAj  )��}�(h�h�j  ]�j  K3j  KAubKBj  )��}�(h�h�j  ]�j  K3j  KBubKCj  )��}�(h�h�j  ]�j  K3j  KCubKDj  )��}�(h�h�j  ]�j  K3j  KDubKEj  )��}�(h�h�j  ]�j  K3j  KEubKFj  )��}�(h�h�j  ]�j  K3j  KFubKGj  )��}�(h�h�j  ]�j  K3j  KGubKHj  )��}�(h�h�j  ]�j  K3j  KHubKIj  )��}�(h�h�j  ]�j  K3j  KIubKJj  )��}�(h�h�j  ]�j  K3j  KJubKKj  )��}�(h�h�j  ]�j  K3j  KKubKLj  )��}�(h�h�j  ]�j  K3j  KLubKMj  )��}�(h�h�j  ]�j  K3j  KMubKNj  )��}�(h�h�j  ]�j  K3j  KNubKOj  )��}�(h�h�j  ]�j  K3j  KOubuK4}�(K j  )��}�(h�h�j  ]�j  K4j  K ubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubK	j  )��}�(h�h�j  ]�j  K4j  K	ubK
j  )��}�(h�h�j  ]�j  K4j  K
ubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�K9aj  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubKj  )��}�(h�h�j  ]�j  K4j  KubK j  )��}�(h�h�j  ]�j  K4j  K ubK!j  )��}�(h�h�j  ]�j  K4j  K!ubK"j  )��}�(h�h�j  ]�j  K4j  K"ubK#j  )��}�(h�h�j  ]�j  K4j  K#ubK$j  )��}�(h�h�j  ]�j  K4j  K$ubK%j  )��}�(h�h�j  ]�j  K4j  K%ubK&j  )��}�(h�h�j  ]�j  K4j  K&ubK'j  )��}�(h�h�j  ]�j  K4j  K'ubK(j  )��}�(h�h�j  ]�j  K4j  K(ubK)j  )��}�(h�h�j  ]�j  K4j  K)ubK*j  )��}�(h�h�j  ]�j  K4j  K*ubK+j  )��}�(h�h�j  ]�j  K4j  K+ubK,j  )��}�(h�h�j  ]�j  K4j  K,ubK-j  )��}�(h�h�j  ]�j  K4j  K-ubK.j  )��}�(h�h�j  ]�j  K4j  K.ubK/j  )��}�(h�h�j  ]�j  K4j  K/ubK0j  )��}�(h�h�j  ]�j  K4j  K0ubK1j  )��}�(h�h�j  ]�j  K4j  K1ubK2j  )��}�(h�h�j  ]�j  K4j  K2ubK3j  )��}�(h�h�j  ]�j  K4j  K3ubK4j  )��}�(h�h�j  ]�j  K4j  K4ubK5j  )��}�(h�h�j  ]�j  K4j  K5ubK6j  )��}�(h�h�j  ]�j  K4j  K6ubK7j  )��}�(h�h�j  ]�j  K4j  K7ubK8j  )��}�(h�h�j  ]�j  K4j  K8ubK9j  )��}�(h�h�j  ]�j  K4j  K9ubK:j  )��}�(h�h�j  ]�j  K4j  K:ubK;j  )��}�(h�h�j  ]�j  K4j  K;ubK<j  )��}�(h�h�j  ]�j  K4j  K<ubK=j  )��}�(h�h�j  ]�j  K4j  K=ubK>j  )��}�(h�h�j  ]�j  K4j  K>ubK?j  )��}�(h�h�j  ]�j  K4j  K?ubK@j  )��}�(h�h�j  ]�j  K4j  K@ubKAj  )��}�(h�h�j  ]�j  K4j  KAubKBj  )��}�(h�h�j  ]�j  K4j  KBubKCj  )��}�(h�h�j  ]�j  K4j  KCubKDj  )��}�(h�h�j  ]�j  K4j  KDubKEj  )��}�(h�h�j  ]�j  K4j  KEubKFj  )��}�(h�h�j  ]�j  K4j  KFubKGj  )��}�(h�h�j  ]�j  K4j  KGubKHj  )��}�(h�h�j  ]�j  K4j  KHubKIj  )��}�(h�h�j  ]�j  K4j  KIubKJj  )��}�(h�h�j  ]�j  K4j  KJubKKj  )��}�(h�h�j  ]�j  K4j  KKubKLj  )��}�(h�h�j  ]�j  K4j  KLubKMj  )��}�(h�h�j  ]�j  K4j  KMubKNj  )��}�(h�h�j  ]�j  K4j  KNubKOj  )��}�(h�h�j  ]�j  K4j  KOubuK5}�(K j  )��}�(h�h�j  ]�j  K5j  K ubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubK	j  )��}�(h�h�j  ]�K:aj  K5j  K	ubK
j  )��}�(h�h�j  ]�K;aj  K5j  K
ubKj  )��}�(h�h�j  ]�K<aj  K5j  KubKj  )��}�(h�h�j  ]�K=aj  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubKj  )��}�(h�h�j  ]�j  K5j  KubK j  )��}�(h�h�j  ]�j  K5j  K ubK!j  )��}�(h�h�j  ]�j  K5j  K!ubK"j  )��}�(h�h�j  ]�j  K5j  K"ubK#j  )��}�(h�h�j  ]�j  K5j  K#ubK$j  )��}�(h�h�j  ]�j  K5j  K$ubK%j  )��}�(h�h�j  ]�j  K5j  K%ubK&j  )��}�(h�h�j  ]�j  K5j  K&ubK'j  )��}�(h�h�j  ]�j  K5j  K'ubK(j  )��}�(h�h�j  ]�j  K5j  K(ubK)j  )��}�(h�h�j  ]�j  K5j  K)ubK*j  )��}�(h�h�j  ]�j  K5j  K*ubK+j  )��}�(h�h�j  ]�j  K5j  K+ubK,j  )��}�(h�h�j  ]�j  K5j  K,ubK-j  )��}�(h�h�j  ]�j  K5j  K-ubK.j  )��}�(h�h�j  ]�j  K5j  K.ubK/j  )��}�(h�h�j  ]�j  K5j  K/ubK0j  )��}�(h�h�j  ]�j  K5j  K0ubK1j  )��}�(h�h�j  ]�j  K5j  K1ubK2j  )��}�(h�h�j  ]�j  K5j  K2ubK3j  )��}�(h�h�j  ]�j  K5j  K3ubK4j  )��}�(h�h�j  ]�j  K5j  K4ubK5j  )��}�(h�h�j  ]�j  K5j  K5ubK6j  )��}�(h�h�j  ]�j  K5j  K6ubK7j  )��}�(h�h�j  ]�j  K5j  K7ubK8j  )��}�(h�h�j  ]�j  K5j  K8ubK9j  )��}�(h�h�j  ]�j  K5j  K9ubK:j  )��}�(h�h�j  ]�j  K5j  K:ubK;j  )��}�(h�h�j  ]�j  K5j  K;ubK<j  )��}�(h�h�j  ]�j  K5j  K<ubK=j  )��}�(h�h�j  ]�j  K5j  K=ubK>j  )��}�(h�h�j  ]�j  K5j  K>ubK?j  )��}�(h�h�j  ]�j  K5j  K?ubK@j  )��}�(h�h�j  ]�j  K5j  K@ubKAj  )��}�(h�h�j  ]�j  K5j  KAubKBj  )��}�(h�h�j  ]�j  K5j  KBubKCj  )��}�(h�h�j  ]�j  K5j  KCubKDj  )��}�(h�h�j  ]�j  K5j  KDubKEj  )��}�(h�h�j  ]�j  K5j  KEubKFj  )��}�(h�h�j  ]�j  K5j  KFubKGj  )��}�(h�h�j  ]�j  K5j  KGubKHj  )��}�(h�h�j  ]�j  K5j  KHubKIj  )��}�(h�h�j  ]�j  K5j  KIubKJj  )��}�(h�h�j  ]�j  K5j  KJubKKj  )��}�(h�h�j  ]�j  K5j  KKubKLj  )��}�(h�h�j  ]�j  K5j  KLubKMj  )��}�(h�h�j  ]�j  K5j  KMubKNj  )��}�(h�h�j  ]�j  K5j  KNubKOj  )��}�(h�h�j  ]�j  K5j  KOubuK6}�(K j  )��}�(h�h�j  ]�j  K6j  K ubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubK	j  )��}�(h�h�j  ]�K>aj  K6j  K	ubK
j  )��}�(h�h�j  ]�j  K6j  K
ubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubKj  )��}�(h�h�j  ]�j  K6j  KubK j  )��}�(h�h�j  ]�j  K6j  K ubK!j  )��}�(h�h�j  ]�j  K6j  K!ubK"j  )��}�(h�h�j  ]�j  K6j  K"ubK#j  )��}�(h�h�j  ]�j  K6j  K#ubK$j  )��}�(h�h�j  ]�j  K6j  K$ubK%j  )��}�(h�h�j  ]�j  K6j  K%ubK&j  )��}�(h�h�j  ]�j  K6j  K&ubK'j  )��}�(h�h�j  ]�j  K6j  K'ubK(j  )��}�(h�h�j  ]�j  K6j  K(ubK)j  )��}�(h�h�j  ]�j  K6j  K)ubK*j  )��}�(h�h�j  ]�j  K6j  K*ubK+j  )��}�(h�h�j  ]�j  K6j  K+ubK,j  )��}�(h�h�j  ]�j  K6j  K,ubK-j  )��}�(h�h�j  ]�j  K6j  K-ubK.j  )��}�(h�h�j  ]�j  K6j  K.ubK/j  )��}�(h�h�j  ]�j  K6j  K/ubK0j  )��}�(h�h�j  ]�j  K6j  K0ubK1j  )��}�(h�h�j  ]�j  K6j  K1ubK2j  )��}�(h�h�j  ]�j  K6j  K2ubK3j  )��}�(h�h�j  ]�j  K6j  K3ubK4j  )��}�(h�h�j  ]�j  K6j  K4ubK5j  )��}�(h�h�j  ]�j  K6j  K5ubK6j  )��}�(h�h�j  ]�j  K6j  K6ubK7j  )��}�(h�h�j  ]�j  K6j  K7ubK8j  )��}�(h�h�j  ]�j  K6j  K8ubK9j  )��}�(h�h�j  ]�j  K6j  K9ubK:j  )��}�(h�h�j  ]�j  K6j  K:ubK;j  )��}�(h�h�j  ]�j  K6j  K;ubK<j  )��}�(h�h�j  ]�j  K6j  K<ubK=j  )��}�(h�h�j  ]�j  K6j  K=ubK>j  )��}�(h�h�j  ]�j  K6j  K>ubK?j  )��}�(h�h�j  ]�j  K6j  K?ubK@j  )��}�(h�h�j  ]�j  K6j  K@ubKAj  )��}�(h�h�j  ]�j  K6j  KAubKBj  )��}�(h�h�j  ]�j  K6j  KBubKCj  )��}�(h�h�j  ]�j  K6j  KCubKDj  )��}�(h�h�j  ]�j  K6j  KDubKEj  )��}�(h�h�j  ]�j  K6j  KEubKFj  )��}�(h�h�j  ]�j  K6j  KFubKGj  )��}�(h�h�j  ]�j  K6j  KGubKHj  )��}�(h�h�j  ]�j  K6j  KHubKIj  )��}�(h�h�j  ]�j  K6j  KIubKJj  )��}�(h�h�j  ]�j  K6j  KJubKKj  )��}�(h�h�j  ]�j  K6j  KKubKLj  )��}�(h�h�j  ]�j  K6j  KLubKMj  )��}�(h�h�j  ]�j  K6j  KMubKNj  )��}�(h�h�j  ]�j  K6j  KNubKOj  )��}�(h�h�j  ]�j  K6j  KOubuK7}�(K j  )��}�(h�h�j  ]�j  K7j  K ubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubK	j  )��}�(h�h�j  ]�j  K7j  K	ubK
j  )��}�(h�h�j  ]�j  K7j  K
ubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubKj  )��}�(h�h�j  ]�j  K7j  KubK j  )��}�(h�h�j  ]�j  K7j  K ubK!j  )��}�(h�h�j  ]�j  K7j  K!ubK"j  )��}�(h�h�j  ]�j  K7j  K"ubK#j  )��}�(h�h�j  ]�j  K7j  K#ubK$j  )��}�(h�h�j  ]�j  K7j  K$ubK%j  )��}�(h�h�j  ]�j  K7j  K%ubK&j  )��}�(h�h�j  ]�j  K7j  K&ubK'j  )��}�(h�h�j  ]�j  K7j  K'ubK(j  )��}�(h�h�j  ]�j  K7j  K(ubK)j  )��}�(h�h�j  ]�j  K7j  K)ubK*j  )��}�(h�h�j  ]�j  K7j  K*ubK+j  )��}�(h�h�j  ]�j  K7j  K+ubK,j  )��}�(h�h�j  ]�j  K7j  K,ubK-j  )��}�(h�h�j  ]�j  K7j  K-ubK.j  )��}�(h�h�j  ]�j  K7j  K.ubK/j  )��}�(h�h�j  ]�j  K7j  K/ubK0j  )��}�(h�h�j  ]�j  K7j  K0ubK1j  )��}�(h�h�j  ]�j  K7j  K1ubK2j  )��}�(h�h�j  ]�j  K7j  K2ubK3j  )��}�(h�h�j  ]�j  K7j  K3ubK4j  )��}�(h�h�j  ]�j  K7j  K4ubK5j  )��}�(h�h�j  ]�j  K7j  K5ubK6j  )��}�(h�h�j  ]�j  K7j  K6ubK7j  )��}�(h�h�j  ]�j  K7j  K7ubK8j  )��}�(h�h�j  ]�j  K7j  K8ubK9j  )��}�(h�h�j  ]�j  K7j  K9ubK:j  )��}�(h�h�j  ]�j  K7j  K:ubK;j  )��}�(h�h�j  ]�j  K7j  K;ubK<j  )��}�(h�h�j  ]�j  K7j  K<ubK=j  )��}�(h�h�j  ]�j  K7j  K=ubK>j  )��}�(h�h�j  ]�j  K7j  K>ubK?j  )��}�(h�h�j  ]�j  K7j  K?ubK@j  )��}�(h�h�j  ]�j  K7j  K@ubKAj  )��}�(h�h�j  ]�j  K7j  KAubKBj  )��}�(h�h�j  ]�j  K7j  KBubKCj  )��}�(h�h�j  ]�j  K7j  KCubKDj  )��}�(h�h�j  ]�j  K7j  KDubKEj  )��}�(h�h�j  ]�j  K7j  KEubKFj  )��}�(h�h�j  ]�j  K7j  KFubKGj  )��}�(h�h�j  ]�j  K7j  KGubKHj  )��}�(h�h�j  ]�j  K7j  KHubKIj  )��}�(h�h�j  ]�j  K7j  KIubKJj  )��}�(h�h�j  ]�j  K7j  KJubKKj  )��}�(h�h�j  ]�j  K7j  KKubKLj  )��}�(h�h�j  ]�j  K7j  KLubKMj  )��}�(h�h�j  ]�j  K7j  KMubKNj  )��}�(h�h�j  ]�j  K7j  KNubKOj  )��}�(h�h�j  ]�j  K7j  KOubuK8}�(K j  )��}�(h�h�j  ]�j  K8j  K ubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubK	j  )��}�(h�h�j  ]�j  K8j  K	ubK
j  )��}�(h�h�j  ]�j  K8j  K
ubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubKj  )��}�(h�h�j  ]�j  K8j  KubK j  )��}�(h�h�j  ]�j  K8j  K ubK!j  )��}�(h�h�j  ]�j  K8j  K!ubK"j  )��}�(h�h�j  ]�j  K8j  K"ubK#j  )��}�(h�h�j  ]�j  K8j  K#ubK$j  )��}�(h�h�j  ]�j  K8j  K$ubK%j  )��}�(h�h�j  ]�j  K8j  K%ubK&j  )��}�(h�h�j  ]�j  K8j  K&ubK'j  )��}�(h�h�j  ]�j  K8j  K'ubK(j  )��}�(h�h�j  ]�j  K8j  K(ubK)j  )��}�(h�h�j  ]�j  K8j  K)ubK*j  )��}�(h�h�j  ]�j  K8j  K*ubK+j  )��}�(h�h�j  ]�j  K8j  K+ubK,j  )��}�(h�h�j  ]�j  K8j  K,ubK-j  )��}�(h�h�j  ]�j  K8j  K-ubK.j  )��}�(h�h�j  ]�j  K8j  K.ubK/j  )��}�(h�h�j  ]�j  K8j  K/ubK0j  )��}�(h�h�j  ]�j  K8j  K0ubK1j  )��}�(h�h�j  ]�j  K8j  K1ubK2j  )��}�(h�h�j  ]�j  K8j  K2ubK3j  )��}�(h�h�j  ]�j  K8j  K3ubK4j  )��}�(h�h�j  ]�j  K8j  K4ubK5j  )��}�(h�h�j  ]�j  K8j  K5ubK6j  )��}�(h�h�j  ]�j  K8j  K6ubK7j  )��}�(h�h�j  ]�j  K8j  K7ubK8j  )��}�(h�h�j  ]�j  K8j  K8ubK9j  )��}�(h�h�j  ]�j  K8j  K9ubK:j  )��}�(h�h�j  ]�j  K8j  K:ubK;j  )��}�(h�h�j  ]�j  K8j  K;ubK<j  )��}�(h�h�j  ]�j  K8j  K<ubK=j  )��}�(h�h�j  ]�j  K8j  K=ubK>j  )��}�(h�h�j  ]�j  K8j  K>ubK?j  )��}�(h�h�j  ]�j  K8j  K?ubK@j  )��}�(h�h�j  ]�j  K8j  K@ubKAj  )��}�(h�h�j  ]�j  K8j  KAubKBj  )��}�(h�h�j  ]�j  K8j  KBubKCj  )��}�(h�h�j  ]�j  K8j  KCubKDj  )��}�(h�h�j  ]�j  K8j  KDubKEj  )��}�(h�h�j  ]�j  K8j  KEubKFj  )��}�(h�h�j  ]�j  K8j  KFubKGj  )��}�(h�h�j  ]�j  K8j  KGubKHj  )��}�(h�h�j  ]�j  K8j  KHubKIj  )��}�(h�h�j  ]�j  K8j  KIubKJj  )��}�(h�h�j  ]�j  K8j  KJubKKj  )��}�(h�h�j  ]�j  K8j  KKubKLj  )��}�(h�h�j  ]�j  K8j  KLubKMj  )��}�(h�h�j  ]�j  K8j  KMubKNj  )��}�(h�h�j  ]�j  K8j  KNubKOj  )��}�(h�h�j  ]�j  K8j  KOubuK9}�(K j  )��}�(h�h�j  ]�j  K9j  K ubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubK	j  )��}�(h�h�j  ]�j  K9j  K	ubK
j  )��}�(h�h�j  ]�j  K9j  K
ubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubKj  )��}�(h�h�j  ]�j  K9j  KubK j  )��}�(h�h�j  ]�j  K9j  K ubK!j  )��}�(h�h�j  ]�j  K9j  K!ubK"j  )��}�(h�h�j  ]�j  K9j  K"ubK#j  )��}�(h�h�j  ]�j  K9j  K#ubK$j  )��}�(h�h�j  ]�j  K9j  K$ubK%j  )��}�(h�h�j  ]�j  K9j  K%ubK&j  )��}�(h�h�j  ]�j  K9j  K&ubK'j  )��}�(h�h�j  ]�j  K9j  K'ubK(j  )��}�(h�h�j  ]�j  K9j  K(ubK)j  )��}�(h�h�j  ]�j  K9j  K)ubK*j  )��}�(h�h�j  ]�j  K9j  K*ubK+j  )��}�(h�h�j  ]�j  K9j  K+ubK,j  )��}�(h�h�j  ]�j  K9j  K,ubK-j  )��}�(h�h�j  ]�j  K9j  K-ubK.j  )��}�(h�h�j  ]�j  K9j  K.ubK/j  )��}�(h�h�j  ]�j  K9j  K/ubK0j  )��}�(h�h�j  ]�j  K9j  K0ubK1j  )��}�(h�h�j  ]�j  K9j  K1ubK2j  )��}�(h�h�j  ]�j  K9j  K2ubK3j  )��}�(h�h�j  ]�j  K9j  K3ubK4j  )��}�(h�h�j  ]�j  K9j  K4ubK5j  )��}�(h�h�j  ]�j  K9j  K5ubK6j  )��}�(h�h�j  ]�j  K9j  K6ubK7j  )��}�(h�h�j  ]�j  K9j  K7ubK8j  )��}�(h�h�j  ]�j  K9j  K8ubK9j  )��}�(h�h�j  ]�j  K9j  K9ubK:j  )��}�(h�h�j  ]�j  K9j  K:ubK;j  )��}�(h�h�j  ]�j  K9j  K;ubK<j  )��}�(h�h�j  ]�j  K9j  K<ubK=j  )��}�(h�h�j  ]�j  K9j  K=ubK>j  )��}�(h�h�j  ]�j  K9j  K>ubK?j  )��}�(h�h�j  ]�j  K9j  K?ubK@j  )��}�(h�h�j  ]�j  K9j  K@ubKAj  )��}�(h�h�j  ]�j  K9j  KAubKBj  )��}�(h�h�j  ]�j  K9j  KBubKCj  )��}�(h�h�j  ]�j  K9j  KCubKDj  )��}�(h�h�j  ]�j  K9j  KDubKEj  )��}�(h�h�j  ]�j  K9j  KEubKFj  )��}�(h�h�j  ]�j  K9j  KFubKGj  )��}�(h�h�j  ]�j  K9j  KGubKHj  )��}�(h�h�j  ]�j  K9j  KHubKIj  )��}�(h�h�j  ]�j  K9j  KIubKJj  )��}�(h�h�j  ]�j  K9j  KJubKKj  )��}�(h�h�j  ]�j  K9j  KKubKLj  )��}�(h�h�j  ]�j  K9j  KLubKMj  )��}�(h�h�j  ]�j  K9j  KMubKNj  )��}�(h�h�j  ]�j  K9j  KNubKOj  )��}�(h�h�j  ]�j  K9j  KOubuK:}�(K j  )��}�(h�h�j  ]�j  K:j  K ubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubK	j  )��}�(h�h�j  ]�j  K:j  K	ubK
j  )��}�(h�h�j  ]�j  K:j  K
ubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubKj  )��}�(h�h�j  ]�j  K:j  KubK j  )��}�(h�h�j  ]�j  K:j  K ubK!j  )��}�(h�h�j  ]�j  K:j  K!ubK"j  )��}�(h�h�j  ]�j  K:j  K"ubK#j  )��}�(h�h�j  ]�j  K:j  K#ubK$j  )��}�(h�h�j  ]�j  K:j  K$ubK%j  )��}�(h�h�j  ]�j  K:j  K%ubK&j  )��}�(h�h�j  ]�j  K:j  K&ubK'j  )��}�(h�h�j  ]�j  K:j  K'ubK(j  )��}�(h�h�j  ]�j  K:j  K(ubK)j  )��}�(h�h�j  ]�j  K:j  K)ubK*j  )��}�(h�h�j  ]�j  K:j  K*ubK+j  )��}�(h�h�j  ]�j  K:j  K+ubK,j  )��}�(h�h�j  ]�j  K:j  K,ubK-j  )��}�(h�h�j  ]�j  K:j  K-ubK.j  )��}�(h�h�j  ]�j  K:j  K.ubK/j  )��}�(h�h�j  ]�j  K:j  K/ubK0j  )��}�(h�h�j  ]�j  K:j  K0ubK1j  )��}�(h�h�j  ]�j  K:j  K1ubK2j  )��}�(h�h�j  ]�j  K:j  K2ubK3j  )��}�(h�h�j  ]�j  K:j  K3ubK4j  )��}�(h�h�j  ]�j  K:j  K4ubK5j  )��}�(h�h�j  ]�j  K:j  K5ubK6j  )��}�(h�h�j  ]�j  K:j  K6ubK7j  )��}�(h�h�j  ]�j  K:j  K7ubK8j  )��}�(h�h�j  ]�j  K:j  K8ubK9j  )��}�(h�h�j  ]�j  K:j  K9ubK:j  )��}�(h�h�j  ]�j  K:j  K:ubK;j  )��}�(h�h�j  ]�j  K:j  K;ubK<j  )��}�(h�h�j  ]�j  K:j  K<ubK=j  )��}�(h�h�j  ]�j  K:j  K=ubK>j  )��}�(h�h�j  ]�j  K:j  K>ubK?j  )��}�(h�h�j  ]�j  K:j  K?ubK@j  )��}�(h�h�j  ]�j  K:j  K@ubKAj  )��}�(h�h�j  ]�j  K:j  KAubKBj  )��}�(h�h�j  ]�j  K:j  KBubKCj  )��}�(h�h�j  ]�j  K:j  KCubKDj  )��}�(h�h�j  ]�j  K:j  KDubKEj  )��}�(h�h�j  ]�j  K:j  KEubKFj  )��}�(h�h�j  ]�j  K:j  KFubKGj  )��}�(h�h�j  ]�j  K:j  KGubKHj  )��}�(h�h�j  ]�j  K:j  KHubKIj  )��}�(h�h�j  ]�j  K:j  KIubKJj  )��}�(h�h�j  ]�j  K:j  KJubKKj  )��}�(h�h�j  ]�j  K:j  KKubKLj  )��}�(h�h�j  ]�j  K:j  KLubKMj  )��}�(h�h�j  ]�j  K:j  KMubKNj  )��}�(h�h�j  ]�j  K:j  KNubKOj  )��}�(h�h�j  ]�j  K:j  KOubuK;}�(K j  )��}�(h�h�j  ]�j  K;j  K ubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubK	j  )��}�(h�h�j  ]�j  K;j  K	ubK
j  )��}�(h�h�j  ]�j  K;j  K
ubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubKj  )��}�(h�h�j  ]�j  K;j  KubK j  )��}�(h�h�j  ]�j  K;j  K ubK!j  )��}�(h�h�j  ]�j  K;j  K!ubK"j  )��}�(h�h�j  ]�j  K;j  K"ubK#j  )��}�(h�h�j  ]�j  K;j  K#ubK$j  )��}�(h�h�j  ]�j  K;j  K$ubK%j  )��}�(h�h�j  ]�j  K;j  K%ubK&j  )��}�(h�h�j  ]�j  K;j  K&ubK'j  )��}�(h�h�j  ]�j  K;j  K'ubK(j  )��}�(h�h�j  ]�j  K;j  K(ubK)j  )��}�(h�h�j  ]�j  K;j  K)ubK*j  )��}�(h�h�j  ]�j  K;j  K*ubK+j  )��}�(h�h�j  ]�j  K;j  K+ubK,j  )��}�(h�h�j  ]�j  K;j  K,ubK-j  )��}�(h�h�j  ]�j  K;j  K-ubK.j  )��}�(h�h�j  ]�j  K;j  K.ubK/j  )��}�(h�h�j  ]�j  K;j  K/ubK0j  )��}�(h�h�j  ]�j  K;j  K0ubK1j  )��}�(h�h�j  ]�j  K;j  K1ubK2j  )��}�(h�h�j  ]�j  K;j  K2ubK3j  )��}�(h�h�j  ]�j  K;j  K3ubK4j  )��}�(h�h�j  ]�j  K;j  K4ubK5j  )��}�(h�h�j  ]�j  K;j  K5ubK6j  )��}�(h�h�j  ]�j  K;j  K6ubK7j  )��}�(h�h�j  ]�j  K;j  K7ubK8j  )��}�(h�h�j  ]�j  K;j  K8ubK9j  )��}�(h�h�j  ]�j  K;j  K9ubK:j  )��}�(h�h�j  ]�j  K;j  K:ubK;j  )��}�(h�h�j  ]�j  K;j  K;ubK<j  )��}�(h�h�j  ]�j  K;j  K<ubK=j  )��}�(h�h�j  ]�j  K;j  K=ubK>j  )��}�(h�h�j  ]�j  K;j  K>ubK?j  )��}�(h�h�j  ]�j  K;j  K?ubK@j  )��}�(h�h�j  ]�j  K;j  K@ubKAj  )��}�(h�h�j  ]�j  K;j  KAubKBj  )��}�(h�h�j  ]�j  K;j  KBubKCj  )��}�(h�h�j  ]�j  K;j  KCubKDj  )��}�(h�h�j  ]�j  K;j  KDubKEj  )��}�(h�h�j  ]�j  K;j  KEubKFj  )��}�(h�h�j  ]�j  K;j  KFubKGj  )��}�(h�h�j  ]�j  K;j  KGubKHj  )��}�(h�h�j  ]�j  K;j  KHubKIj  )��}�(h�h�j  ]�j  K;j  KIubKJj  )��}�(h�h�j  ]�j  K;j  KJubKKj  )��}�(h�h�j  ]�j  K;j  KKubKLj  )��}�(h�h�j  ]�j  K;j  KLubKMj  )��}�(h�h�j  ]�j  K;j  KMubKNj  )��}�(h�h�j  ]�j  K;j  KNubKOj  )��}�(h�h�j  ]�j  K;j  KOubuK<}�(K j  )��}�(h�h�j  ]�j  K<j  K ubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubK	j  )��}�(h�h�j  ]�j  K<j  K	ubK
j  )��}�(h�h�j  ]�j  K<j  K
ubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubKj  )��}�(h�h�j  ]�j  K<j  KubK j  )��}�(h�h�j  ]�j  K<j  K ubK!j  )��}�(h�h�j  ]�j  K<j  K!ubK"j  )��}�(h�h�j  ]�j  K<j  K"ubK#j  )��}�(h�h�j  ]�j  K<j  K#ubK$j  )��}�(h�h�j  ]�j  K<j  K$ubK%j  )��}�(h�h�j  ]�j  K<j  K%ubK&j  )��}�(h�h�j  ]�j  K<j  K&ubK'j  )��}�(h�h�j  ]�j  K<j  K'ubK(j  )��}�(h�h�j  ]�j  K<j  K(ubK)j  )��}�(h�h�j  ]�j  K<j  K)ubK*j  )��}�(h�h�j  ]�j  K<j  K*ubK+j  )��}�(h�h�j  ]�j  K<j  K+ubK,j  )��}�(h�h�j  ]�j  K<j  K,ubK-j  )��}�(h�h�j  ]�j  K<j  K-ubK.j  )��}�(h�h�j  ]�j  K<j  K.ubK/j  )��}�(h�h�j  ]�j  K<j  K/ubK0j  )��}�(h�h�j  ]�j  K<j  K0ubK1j  )��}�(h�h�j  ]�j  K<j  K1ubK2j  )��}�(h�h�j  ]�j  K<j  K2ubK3j  )��}�(h�h�j  ]�j  K<j  K3ubK4j  )��}�(h�h�j  ]�j  K<j  K4ubK5j  )��}�(h�h�j  ]�j  K<j  K5ubK6j  )��}�(h�h�j  ]�j  K<j  K6ubK7j  )��}�(h�h�j  ]�j  K<j  K7ubK8j  )��}�(h�h�j  ]�j  K<j  K8ubK9j  )��}�(h�h�j  ]�j  K<j  K9ubK:j  )��}�(h�h�j  ]�j  K<j  K:ubK;j  )��}�(h�h�j  ]�j  K<j  K;ubK<j  )��}�(h�h�j  ]�j  K<j  K<ubK=j  )��}�(h�h�j  ]�j  K<j  K=ubK>j  )��}�(h�h�j  ]�j  K<j  K>ubK?j  )��}�(h�h�j  ]�j  K<j  K?ubK@j  )��}�(h�h�j  ]�j  K<j  K@ubKAj  )��}�(h�h�j  ]�j  K<j  KAubKBj  )��}�(h�h�j  ]�j  K<j  KBubKCj  )��}�(h�h�j  ]�j  K<j  KCubKDj  )��}�(h�h�j  ]�j  K<j  KDubKEj  )��}�(h�h�j  ]�j  K<j  KEubKFj  )��}�(h�h�j  ]�j  K<j  KFubKGj  )��}�(h�h�j  ]�j  K<j  KGubKHj  )��}�(h�h�j  ]�j  K<j  KHubKIj  )��}�(h�h�j  ]�j  K<j  KIubKJj  )��}�(h�h�j  ]�j  K<j  KJubKKj  )��}�(h�h�j  ]�j  K<j  KKubKLj  )��}�(h�h�j  ]�j  K<j  KLubKMj  )��}�(h�h�j  ]�j  K<j  KMubKNj  )��}�(h�h�j  ]�j  K<j  KNubKOj  )��}�(h�h�j  ]�j  K<j  KOubuK=}�(K j  )��}�(h�h�j  ]�j  K=j  K ubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubK	j  )��}�(h�h�j  ]�K?aj  K=j  K	ubK
j  )��}�(h�h�j  ]�j  K=j  K
ubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubKj  )��}�(h�h�j  ]�j  K=j  KubK j  )��}�(h�h�j  ]�j  K=j  K ubK!j  )��}�(h�h�j  ]�j  K=j  K!ubK"j  )��}�(h�h�j  ]�j  K=j  K"ubK#j  )��}�(h�h�j  ]�j  K=j  K#ubK$j  )��}�(h�h�j  ]�j  K=j  K$ubK%j  )��}�(h�h�j  ]�j  K=j  K%ubK&j  )��}�(h�h�j  ]�j  K=j  K&ubK'j  )��}�(h�h�j  ]�j  K=j  K'ubK(j  )��}�(h�h�j  ]�j  K=j  K(ubK)j  )��}�(h�h�j  ]�j  K=j  K)ubK*j  )��}�(h�h�j  ]�j  K=j  K*ubK+j  )��}�(h�h�j  ]�j  K=j  K+ubK,j  )��}�(h�h�j  ]�j  K=j  K,ubK-j  )��}�(h�h�j  ]�j  K=j  K-ubK.j  )��}�(h�h�j  ]�j  K=j  K.ubK/j  )��}�(h�h�j  ]�j  K=j  K/ubK0j  )��}�(h�h�j  ]�j  K=j  K0ubK1j  )��}�(h�h�j  ]�j  K=j  K1ubK2j  )��}�(h�h�j  ]�j  K=j  K2ubK3j  )��}�(h�h�j  ]�j  K=j  K3ubK4j  )��}�(h�h�j  ]�j  K=j  K4ubK5j  )��}�(h�h�j  ]�j  K=j  K5ubK6j  )��}�(h�h�j  ]�j  K=j  K6ubK7j  )��}�(h�h�j  ]�j  K=j  K7ubK8j  )��}�(h�h�j  ]�j  K=j  K8ubK9j  )��}�(h�h�j  ]�j  K=j  K9ubK:j  )��}�(h�h�j  ]�j  K=j  K:ubK;j  )��}�(h�h�j  ]�j  K=j  K;ubK<j  )��}�(h�h�j  ]�j  K=j  K<ubK=j  )��}�(h�h�j  ]�j  K=j  K=ubK>j  )��}�(h�h�j  ]�j  K=j  K>ubK?j  )��}�(h�h�j  ]�j  K=j  K?ubK@j  )��}�(h�h�j  ]�j  K=j  K@ubKAj  )��}�(h�h�j  ]�j  K=j  KAubKBj  )��}�(h�h�j  ]�j  K=j  KBubKCj  )��}�(h�h�j  ]�j  K=j  KCubKDj  )��}�(h�h�j  ]�j  K=j  KDubKEj  )��}�(h�h�j  ]�j  K=j  KEubKFj  )��}�(h�h�j  ]�j  K=j  KFubKGj  )��}�(h�h�j  ]�j  K=j  KGubKHj  )��}�(h�h�j  ]�j  K=j  KHubKIj  )��}�(h�h�j  ]�j  K=j  KIubKJj  )��}�(h�h�j  ]�j  K=j  KJubKKj  )��}�(h�h�j  ]�j  K=j  KKubKLj  )��}�(h�h�j  ]�j  K=j  KLubKMj  )��}�(h�h�j  ]�j  K=j  KMubKNj  )��}�(h�h�j  ]�j  K=j  KNubKOj  )��}�(h�h�j  ]�j  K=j  KOubuK>}�(K j  )��}�(h�h�j  ]�j  K>j  K ubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubK	j  )��}�(h�h�j  ]�j  K>j  K	ubK
j  )��}�(h�h�j  ]�K@aj  K>j  K
ubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubKj  )��}�(h�h�j  ]�j  K>j  KubK j  )��}�(h�h�j  ]�j  K>j  K ubK!j  )��}�(h�h�j  ]�j  K>j  K!ubK"j  )��}�(h�h�j  ]�j  K>j  K"ubK#j  )��}�(h�h�j  ]�j  K>j  K#ubK$j  )��}�(h�h�j  ]�j  K>j  K$ubK%j  )��}�(h�h�j  ]�j  K>j  K%ubK&j  )��}�(h�h�j  ]�j  K>j  K&ubK'j  )��}�(h�h�j  ]�j  K>j  K'ubK(j  )��}�(h�h�j  ]�j  K>j  K(ubK)j  )��}�(h�h�j  ]�j  K>j  K)ubK*j  )��}�(h�h�j  ]�j  K>j  K*ubK+j  )��}�(h�h�j  ]�j  K>j  K+ubK,j  )��}�(h�h�j  ]�j  K>j  K,ubK-j  )��}�(h�h�j  ]�j  K>j  K-ubK.j  )��}�(h�h�j  ]�j  K>j  K.ubK/j  )��}�(h�h�j  ]�j  K>j  K/ubK0j  )��}�(h�h�j  ]�j  K>j  K0ubK1j  )��}�(h�h�j  ]�j  K>j  K1ubK2j  )��}�(h�h�j  ]�j  K>j  K2ubK3j  )��}�(h�h�j  ]�j  K>j  K3ubK4j  )��}�(h�h�j  ]�j  K>j  K4ubK5j  )��}�(h�h�j  ]�j  K>j  K5ubK6j  )��}�(h�h�j  ]�j  K>j  K6ubK7j  )��}�(h�h�j  ]�j  K>j  K7ubK8j  )��}�(h�h�j  ]�j  K>j  K8ubK9j  )��}�(h�h�j  ]�j  K>j  K9ubK:j  )��}�(h�h�j  ]�j  K>j  K:ubK;j  )��}�(h�h�j  ]�j  K>j  K;ubK<j  )��}�(h�h�j  ]�j  K>j  K<ubK=j  )��}�(h�h�j  ]�j  K>j  K=ubK>j  )��}�(h�h�j  ]�j  K>j  K>ubK?j  )��}�(h�h�j  ]�j  K>j  K?ubK@j  )��}�(h�h�j  ]�j  K>j  K@ubKAj  )��}�(h�h�j  ]�j  K>j  KAubKBj  )��}�(h�h�j  ]�j  K>j  KBubKCj  )��}�(h�h�j  ]�j  K>j  KCubKDj  )��}�(h�h�j  ]�j  K>j  KDubKEj  )��}�(h�h�j  ]�j  K>j  KEubKFj  )��}�(h�h�j  ]�j  K>j  KFubKGj  )��}�(h�h�j  ]�j  K>j  KGubKHj  )��}�(h�h�j  ]�j  K>j  KHubKIj  )��}�(h�h�j  ]�j  K>j  KIubKJj  )��}�(h�h�j  ]�j  K>j  KJubKKj  )��}�(h�h�j  ]�j  K>j  KKubKLj  )��}�(h�h�j  ]�j  K>j  KLubKMj  )��}�(h�h�j  ]�j  K>j  KMubKNj  )��}�(h�h�j  ]�j  K>j  KNubKOj  )��}�(h�h�j  ]�j  K>j  KOubuK?}�(K j  )��}�(h�h�j  ]�j  K?j  K ubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubK	j  )��}�(h�h�j  ]�KCaj  K?j  K	ubK
j  )��}�(h�h�j  ]�j  K?j  K
ubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubKj  )��}�(h�h�j  ]�j  K?j  KubK j  )��}�(h�h�j  ]�j  K?j  K ubK!j  )��}�(h�h�j  ]�j  K?j  K!ubK"j  )��}�(h�h�j  ]�j  K?j  K"ubK#j  )��}�(h�h�j  ]�j  K?j  K#ubK$j  )��}�(h�h�j  ]�j  K?j  K$ubK%j  )��}�(h�h�j  ]�j  K?j  K%ubK&j  )��}�(h�h�j  ]�j  K?j  K&ubK'j  )��}�(h�h�j  ]�j  K?j  K'ubK(j  )��}�(h�h�j  ]�j  K?j  K(ubK)j  )��}�(h�h�j  ]�j  K?j  K)ubK*j  )��}�(h�h�j  ]�j  K?j  K*ubK+j  )��}�(h�h�j  ]�j  K?j  K+ubK,j  )��}�(h�h�j  ]�j  K?j  K,ubK-j  )��}�(h�h�j  ]�j  K?j  K-ubK.j  )��}�(h�h�j  ]�j  K?j  K.ubK/j  )��}�(h�h�j  ]�j  K?j  K/ubK0j  )��}�(h�h�j  ]�j  K?j  K0ubK1j  )��}�(h�h�j  ]�j  K?j  K1ubK2j  )��}�(h�h�j  ]�j  K?j  K2ubK3j  )��}�(h�h�j  ]�j  K?j  K3ubK4j  )��}�(h�h�j  ]�j  K?j  K4ubK5j  )��}�(h�h�j  ]�j  K?j  K5ubK6j  )��}�(h�h�j  ]�j  K?j  K6ubK7j  )��}�(h�h�j  ]�j  K?j  K7ubK8j  )��}�(h�h�j  ]�j  K?j  K8ubK9j  )��}�(h�h�j  ]�j  K?j  K9ubK:j  )��}�(h�h�j  ]�j  K?j  K:ubK;j  )��}�(h�h�j  ]�j  K?j  K;ubK<j  )��}�(h�h�j  ]�j  K?j  K<ubK=j  )��}�(h�h�j  ]�j  K?j  K=ubK>j  )��}�(h�h�j  ]�j  K?j  K>ubK?j  )��}�(h�h�j  ]�j  K?j  K?ubK@j  )��}�(h�h�j  ]�j  K?j  K@ubKAj  )��}�(h�h�j  ]�j  K?j  KAubKBj  )��}�(h�h�j  ]�j  K?j  KBubKCj  )��}�(h�h�j  ]�j  K?j  KCubKDj  )��}�(h�h�j  ]�j  K?j  KDubKEj  )��}�(h�h�j  ]�j  K?j  KEubKFj  )��}�(h�h�j  ]�j  K?j  KFubKGj  )��}�(h�h�j  ]�j  K?j  KGubKHj  )��}�(h�h�j  ]�j  K?j  KHubKIj  )��}�(h�h�j  ]�j  K?j  KIubKJj  )��}�(h�h�j  ]�j  K?j  KJubKKj  )��}�(h�h�j  ]�j  K?j  KKubKLj  )��}�(h�h�j  ]�j  K?j  KLubKMj  )��}�(h�h�j  ]�j  K?j  KMubKNj  )��}�(h�h�j  ]�j  K?j  KNubKOj  )��}�(h�h�j  ]�j  K?j  KOubuK@}�(K j  )��}�(h�h�j  ]�j  K@j  K ubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubK	j  )��}�(h�h�j  ]�j  K@j  K	ubK
j  )��}�(h�h�j  ]�KDaj  K@j  K
ubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubKj  )��}�(h�h�j  ]�j  K@j  KubK j  )��}�(h�h�j  ]�j  K@j  K ubK!j  )��}�(h�h�j  ]�j  K@j  K!ubK"j  )��}�(h�h�j  ]�j  K@j  K"ubK#j  )��}�(h�h�j  ]�j  K@j  K#ubK$j  )��}�(h�h�j  ]�j  K@j  K$ubK%j  )��}�(h�h�j  ]�j  K@j  K%ubK&j  )��}�(h�h�j  ]�j  K@j  K&ubK'j  )��}�(h�h�j  ]�j  K@j  K'ubK(j  )��}�(h�h�j  ]�j  K@j  K(ubK)j  )��}�(h�h�j  ]�j  K@j  K)ubK*j  )��}�(h�h�j  ]�j  K@j  K*ubK+j  )��}�(h�h�j  ]�j  K@j  K+ubK,j  )��}�(h�h�j  ]�j  K@j  K,ubK-j  )��}�(h�h�j  ]�j  K@j  K-ubK.j  )��}�(h�h�j  ]�j  K@j  K.ubK/j  )��}�(h�h�j  ]�j  K@j  K/ubK0j  )��}�(h�h�j  ]�j  K@j  K0ubK1j  )��}�(h�h�j  ]�j  K@j  K1ubK2j  )��}�(h�h�j  ]�j  K@j  K2ubK3j  )��}�(h�h�j  ]�j  K@j  K3ubK4j  )��}�(h�h�j  ]�j  K@j  K4ubK5j  )��}�(h�h�j  ]�j  K@j  K5ubK6j  )��}�(h�h�j  ]�j  K@j  K6ubK7j  )��}�(h�h�j  ]�j  K@j  K7ubK8j  )��}�(h�h�j  ]�j  K@j  K8ubK9j  )��}�(h�h�j  ]�j  K@j  K9ubK:j  )��}�(h�h�j  ]�j  K@j  K:ubK;j  )��}�(h�h�j  ]�j  K@j  K;ubK<j  )��}�(h�h�j  ]�j  K@j  K<ubK=j  )��}�(h�h�j  ]�j  K@j  K=ubK>j  )��}�(h�h�j  ]�j  K@j  K>ubK?j  )��}�(h�h�j  ]�j  K@j  K?ubK@j  )��}�(h�h�j  ]�j  K@j  K@ubKAj  )��}�(h�h�j  ]�j  K@j  KAubKBj  )��}�(h�h�j  ]�j  K@j  KBubKCj  )��}�(h�h�j  ]�j  K@j  KCubKDj  )��}�(h�h�j  ]�j  K@j  KDubKEj  )��}�(h�h�j  ]�j  K@j  KEubKFj  )��}�(h�h�j  ]�j  K@j  KFubKGj  )��}�(h�h�j  ]�j  K@j  KGubKHj  )��}�(h�h�j  ]�j  K@j  KHubKIj  )��}�(h�h�j  ]�j  K@j  KIubKJj  )��}�(h�h�j  ]�j  K@j  KJubKKj  )��}�(h�h�j  ]�j  K@j  KKubKLj  )��}�(h�h�j  ]�j  K@j  KLubKMj  )��}�(h�h�j  ]�j  K@j  KMubKNj  )��}�(h�h�j  ]�j  K@j  KNubKOj  )��}�(h�h�j  ]�j  K@j  KOubuKA}�(K j  )��}�(h�h�j  ]�j  KAj  K ubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubK	j  )��}�(h�h�j  ]�j  KAj  K	ubK
j  )��}�(h�h�j  ]�j  KAj  K
ubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubKj  )��}�(h�h�j  ]�j  KAj  KubK j  )��}�(h�h�j  ]�j  KAj  K ubK!j  )��}�(h�h�j  ]�j  KAj  K!ubK"j  )��}�(h�h�j  ]�j  KAj  K"ubK#j  )��}�(h�h�j  ]�j  KAj  K#ubK$j  )��}�(h�h�j  ]�j  KAj  K$ubK%j  )��}�(h�h�j  ]�j  KAj  K%ubK&j  )��}�(h�h�j  ]�j  KAj  K&ubK'j  )��}�(h�h�j  ]�j  KAj  K'ubK(j  )��}�(h�h�j  ]�j  KAj  K(ubK)j  )��}�(h�h�j  ]�j  KAj  K)ubK*j  )��}�(h�h�j  ]�j  KAj  K*ubK+j  )��}�(h�h�j  ]�j  KAj  K+ubK,j  )��}�(h�h�j  ]�j  KAj  K,ubK-j  )��}�(h�h�j  ]�j  KAj  K-ubK.j  )��}�(h�h�j  ]�j  KAj  K.ubK/j  )��}�(h�h�j  ]�j  KAj  K/ubK0j  )��}�(h�h�j  ]�j  KAj  K0ubK1j  )��}�(h�h�j  ]�j  KAj  K1ubK2j  )��}�(h�h�j  ]�KEaj  KAj  K2ubK3j  )��}�(h�h�j  ]�j  KAj  K3ubK4j  )��}�(h�h�j  ]�j  KAj  K4ubK5j  )��}�(h�h�j  ]�j  KAj  K5ubK6j  )��}�(h�h�j  ]�j  KAj  K6ubK7j  )��}�(h�h�j  ]�j  KAj  K7ubK8j  )��}�(h�h�j  ]�j  KAj  K8ubK9j  )��}�(h�h�j  ]�j  KAj  K9ubK:j  )��}�(h�h�j  ]�j  KAj  K:ubK;j  )��}�(h�h�j  ]�j  KAj  K;ubK<j  )��}�(h�h�j  ]�j  KAj  K<ubK=j  )��}�(h�h�j  ]�j  KAj  K=ubK>j  )��}�(h�h�j  ]�j  KAj  K>ubK?j  )��}�(h�h�j  ]�j  KAj  K?ubK@j  )��}�(h�h�j  ]�j  KAj  K@ubKAj  )��}�(h�h�j  ]�j  KAj  KAubKBj  )��}�(h�h�j  ]�j  KAj  KBubKCj  )��}�(h�h�j  ]�j  KAj  KCubKDj  )��}�(h�h�j  ]�j  KAj  KDubKEj  )��}�(h�h�j  ]�j  KAj  KEubKFj  )��}�(h�h�j  ]�j  KAj  KFubKGj  )��}�(h�h�j  ]�j  KAj  KGubKHj  )��}�(h�h�j  ]�j  KAj  KHubKIj  )��}�(h�h�j  ]�j  KAj  KIubKJj  )��}�(h�h�j  ]�j  KAj  KJubKKj  )��}�(h�h�j  ]�j  KAj  KKubKLj  )��}�(h�h�j  ]�j  KAj  KLubKMj  )��}�(h�h�j  ]�j  KAj  KMubKNj  )��}�(h�h�j  ]�j  KAj  KNubKOj  )��}�(h�h�j  ]�j  KAj  KOubuKB}�(K j  )��}�(h�h�j  ]�j  KBj  K ubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubK	j  )��}�(h�h�j  ]�j  KBj  K	ubK
j  )��}�(h�h�j  ]�KFaj  KBj  K
ubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubKj  )��}�(h�h�j  ]�j  KBj  KubK j  )��}�(h�h�j  ]�j  KBj  K ubK!j  )��}�(h�h�j  ]�j  KBj  K!ubK"j  )��}�(h�h�j  ]�j  KBj  K"ubK#j  )��}�(h�h�j  ]�j  KBj  K#ubK$j  )��}�(h�h�j  ]�j  KBj  K$ubK%j  )��}�(h�h�j  ]�j  KBj  K%ubK&j  )��}�(h�h�j  ]�j  KBj  K&ubK'j  )��}�(h�h�j  ]�j  KBj  K'ubK(j  )��}�(h�h�j  ]�j  KBj  K(ubK)j  )��}�(h�h�j  ]�j  KBj  K)ubK*j  )��}�(h�h�j  ]�j  KBj  K*ubK+j  )��}�(h�h�j  ]�j  KBj  K+ubK,j  )��}�(h�h�j  ]�j  KBj  K,ubK-j  )��}�(h�h�j  ]�j  KBj  K-ubK.j  )��}�(h�h�j  ]�j  KBj  K.ubK/j  )��}�(h�h�j  ]�j  KBj  K/ubK0j  )��}�(h�h�j  ]�j  KBj  K0ubK1j  )��}�(h�h�j  ]�j  KBj  K1ubK2j  )��}�(h�h�j  ]�j  KBj  K2ubK3j  )��}�(h�h�j  ]�j  KBj  K3ubK4j  )��}�(h�h�j  ]�j  KBj  K4ubK5j  )��}�(h�h�j  ]�j  KBj  K5ubK6j  )��}�(h�h�j  ]�j  KBj  K6ubK7j  )��}�(h�h�j  ]�j  KBj  K7ubK8j  )��}�(h�h�j  ]�j  KBj  K8ubK9j  )��}�(h�h�j  ]�j  KBj  K9ubK:j  )��}�(h�h�j  ]�j  KBj  K:ubK;j  )��}�(h�h�j  ]�j  KBj  K;ubK<j  )��}�(h�h�j  ]�j  KBj  K<ubK=j  )��}�(h�h�j  ]�j  KBj  K=ubK>j  )��}�(h�h�j  ]�j  KBj  K>ubK?j  )��}�(h�h�j  ]�j  KBj  K?ubK@j  )��}�(h�h�j  ]�j  KBj  K@ubKAj  )��}�(h�h�j  ]�j  KBj  KAubKBj  )��}�(h�h�j  ]�j  KBj  KBubKCj  )��}�(h�h�j  ]�j  KBj  KCubKDj  )��}�(h�h�j  ]�j  KBj  KDubKEj  )��}�(h�h�j  ]�j  KBj  KEubKFj  )��}�(h�h�j  ]�j  KBj  KFubKGj  )��}�(h�h�j  ]�j  KBj  KGubKHj  )��}�(h�h�j  ]�j  KBj  KHubKIj  )��}�(h�h�j  ]�j  KBj  KIubKJj  )��}�(h�h�j  ]�j  KBj  KJubKKj  )��}�(h�h�j  ]�j  KBj  KKubKLj  )��}�(h�h�j  ]�j  KBj  KLubKMj  )��}�(h�h�j  ]�j  KBj  KMubKNj  )��}�(h�h�j  ]�j  KBj  KNubKOj  )��}�(h�h�j  ]�j  KBj  KOubuKC}�(K j  )��}�(h�h�j  ]�j  KCj  K ubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubK	j  )��}�(h�h�j  ]�j  KCj  K	ubK
j  )��}�(h�h�j  ]�KGaj  KCj  K
ubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubKj  )��}�(h�h�j  ]�j  KCj  KubK j  )��}�(h�h�j  ]�j  KCj  K ubK!j  )��}�(h�h�j  ]�j  KCj  K!ubK"j  )��}�(h�h�j  ]�j  KCj  K"ubK#j  )��}�(h�h�j  ]�j  KCj  K#ubK$j  )��}�(h�h�j  ]�j  KCj  K$ubK%j  )��}�(h�h�j  ]�j  KCj  K%ubK&j  )��}�(h�h�j  ]�j  KCj  K&ubK'j  )��}�(h�h�j  ]�j  KCj  K'ubK(j  )��}�(h�h�j  ]�j  KCj  K(ubK)j  )��}�(h�h�j  ]�j  KCj  K)ubK*j  )��}�(h�h�j  ]�j  KCj  K*ubK+j  )��}�(h�h�j  ]�j  KCj  K+ubK,j  )��}�(h�h�j  ]�j  KCj  K,ubK-j  )��}�(h�h�j  ]�j  KCj  K-ubK.j  )��}�(h�h�j  ]�j  KCj  K.ubK/j  )��}�(h�h�j  ]�j  KCj  K/ubK0j  )��}�(h�h�j  ]�j  KCj  K0ubK1j  )��}�(h�h�j  ]�j  KCj  K1ubK2j  )��}�(h�h�j  ]�j  KCj  K2ubK3j  )��}�(h�h�j  ]�j  KCj  K3ubK4j  )��}�(h�h�j  ]�j  KCj  K4ubK5j  )��}�(h�h�j  ]�j  KCj  K5ubK6j  )��}�(h�h�j  ]�j  KCj  K6ubK7j  )��}�(h�h�j  ]�j  KCj  K7ubK8j  )��}�(h�h�j  ]�j  KCj  K8ubK9j  )��}�(h�h�j  ]�j  KCj  K9ubK:j  )��}�(h�h�j  ]�j  KCj  K:ubK;j  )��}�(h�h�j  ]�j  KCj  K;ubK<j  )��}�(h�h�j  ]�j  KCj  K<ubK=j  )��}�(h�h�j  ]�j  KCj  K=ubK>j  )��}�(h�h�j  ]�j  KCj  K>ubK?j  )��}�(h�h�j  ]�j  KCj  K?ubK@j  )��}�(h�h�j  ]�j  KCj  K@ubKAj  )��}�(h�h�j  ]�j  KCj  KAubKBj  )��}�(h�h�j  ]�j  KCj  KBubKCj  )��}�(h�h�j  ]�j  KCj  KCubKDj  )��}�(h�h�j  ]�j  KCj  KDubKEj  )��}�(h�h�j  ]�j  KCj  KEubKFj  )��}�(h�h�j  ]�j  KCj  KFubKGj  )��}�(h�h�j  ]�j  KCj  KGubKHj  )��}�(h�h�j  ]�j  KCj  KHubKIj  )��}�(h�h�j  ]�j  KCj  KIubKJj  )��}�(h�h�j  ]�j  KCj  KJubKKj  )��}�(h�h�j  ]�j  KCj  KKubKLj  )��}�(h�h�j  ]�j  KCj  KLubKMj  )��}�(h�h�j  ]�j  KCj  KMubKNj  )��}�(h�h�j  ]�j  KCj  KNubKOj  )��}�(h�h�j  ]�j  KCj  KOubuKD}�(K j  )��}�(h�h�j  ]�j  KDj  K ubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubK	j  )��}�(h�h�j  ]�j  KDj  K	ubK
j  )��}�(h�h�j  ]�j  KDj  K
ubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubKj  )��}�(h�h�j  ]�j  KDj  KubK j  )��}�(h�h�j  ]�j  KDj  K ubK!j  )��}�(h�h�j  ]�j  KDj  K!ubK"j  )��}�(h�h�j  ]�j  KDj  K"ubK#j  )��}�(h�h�j  ]�j  KDj  K#ubK$j  )��}�(h�h�j  ]�j  KDj  K$ubK%j  )��}�(h�h�j  ]�j  KDj  K%ubK&j  )��}�(h�h�j  ]�j  KDj  K&ubK'j  )��}�(h�h�j  ]�j  KDj  K'ubK(j  )��}�(h�h�j  ]�j  KDj  K(ubK)j  )��}�(h�h�j  ]�j  KDj  K)ubK*j  )��}�(h�h�j  ]�j  KDj  K*ubK+j  )��}�(h�h�j  ]�j  KDj  K+ubK,j  )��}�(h�h�j  ]�KHaj  KDj  K,ubK-j  )��}�(h�h�j  ]�j  KDj  K-ubK.j  )��}�(h�h�j  ]�j  KDj  K.ubK/j  )��}�(h�h�j  ]�j  KDj  K/ubK0j  )��}�(h�h�j  ]�j  KDj  K0ubK1j  )��}�(h�h�j  ]�j  KDj  K1ubK2j  )��}�(h�h�j  ]�j  KDj  K2ubK3j  )��}�(h�h�j  ]�j  KDj  K3ubK4j  )��}�(h�h�j  ]�j  KDj  K4ubK5j  )��}�(h�h�j  ]�j  KDj  K5ubK6j  )��}�(h�h�j  ]�j  KDj  K6ubK7j  )��}�(h�h�j  ]�j  KDj  K7ubK8j  )��}�(h�h�j  ]�j  KDj  K8ubK9j  )��}�(h�h�j  ]�j  KDj  K9ubK:j  )��}�(h�h�j  ]�j  KDj  K:ubK;j  )��}�(h�h�j  ]�j  KDj  K;ubK<j  )��}�(h�h�j  ]�j  KDj  K<ubK=j  )��}�(h�h�j  ]�j  KDj  K=ubK>j  )��}�(h�h�j  ]�j  KDj  K>ubK?j  )��}�(h�h�j  ]�j  KDj  K?ubK@j  )��}�(h�h�j  ]�j  KDj  K@ubKAj  )��}�(h�h�j  ]�j  KDj  KAubKBj  )��}�(h�h�j  ]�j  KDj  KBubKCj  )��}�(h�h�j  ]�j  KDj  KCubKDj  )��}�(h�h�j  ]�j  KDj  KDubKEj  )��}�(h�h�j  ]�j  KDj  KEubKFj  )��}�(h�h�j  ]�j  KDj  KFubKGj  )��}�(h�h�j  ]�j  KDj  KGubKHj  )��}�(h�h�j  ]�j  KDj  KHubKIj  )��}�(h�h�j  ]�j  KDj  KIubKJj  )��}�(h�h�j  ]�j  KDj  KJubKKj  )��}�(h�h�j  ]�j  KDj  KKubKLj  )��}�(h�h�j  ]�j  KDj  KLubKMj  )��}�(h�h�j  ]�j  KDj  KMubKNj  )��}�(h�h�j  ]�j  KDj  KNubKOj  )��}�(h�h�j  ]�j  KDj  KOubuKE}�(K j  )��}�(h�h�j  ]�j  KEj  K ubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubK	j  )��}�(h�h�j  ]�j  KEj  K	ubK
j  )��}�(h�h�j  ]�j  KEj  K
ubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�K7aj  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubKj  )��}�(h�h�j  ]�j  KEj  KubK j  )��}�(h�h�j  ]�j  KEj  K ubK!j  )��}�(h�h�j  ]�j  KEj  K!ubK"j  )��}�(h�h�j  ]�j  KEj  K"ubK#j  )��}�(h�h�j  ]�j  KEj  K#ubK$j  )��}�(h�h�j  ]�j  KEj  K$ubK%j  )��}�(h�h�j  ]�j  KEj  K%ubK&j  )��}�(h�h�j  ]�j  KEj  K&ubK'j  )��}�(h�h�j  ]�j  KEj  K'ubK(j  )��}�(h�h�j  ]�j  KEj  K(ubK)j  )��}�(h�h�j  ]�j  KEj  K)ubK*j  )��}�(h�h�j  ]�j  KEj  K*ubK+j  )��}�(h�h�j  ]�j  KEj  K+ubK,j  )��}�(h�h�j  ]�j  KEj  K,ubK-j  )��}�(h�h�j  ]�j  KEj  K-ubK.j  )��}�(h�h�j  ]�j  KEj  K.ubK/j  )��}�(h�h�j  ]�j  KEj  K/ubK0j  )��}�(h�h�j  ]�j  KEj  K0ubK1j  )��}�(h�h�j  ]�j  KEj  K1ubK2j  )��}�(h�h�j  ]�j  KEj  K2ubK3j  )��}�(h�h�j  ]�j  KEj  K3ubK4j  )��}�(h�h�j  ]�j  KEj  K4ubK5j  )��}�(h�h�j  ]�j  KEj  K5ubK6j  )��}�(h�h�j  ]�j  KEj  K6ubK7j  )��}�(h�h�j  ]�j  KEj  K7ubK8j  )��}�(h�h�j  ]�j  KEj  K8ubK9j  )��}�(h�h�j  ]�j  KEj  K9ubK:j  )��}�(h�h�j  ]�j  KEj  K:ubK;j  )��}�(h�h�j  ]�j  KEj  K;ubK<j  )��}�(h�h�j  ]�j  KEj  K<ubK=j  )��}�(h�h�j  ]�j  KEj  K=ubK>j  )��}�(h�h�j  ]�j  KEj  K>ubK?j  )��}�(h�h�j  ]�j  KEj  K?ubK@j  )��}�(h�h�j  ]�j  KEj  K@ubKAj  )��}�(h�h�j  ]�j  KEj  KAubKBj  )��}�(h�h�j  ]�j  KEj  KBubKCj  )��}�(h�h�j  ]�j  KEj  KCubKDj  )��}�(h�h�j  ]�j  KEj  KDubKEj  )��}�(h�h�j  ]�j  KEj  KEubKFj  )��}�(h�h�j  ]�j  KEj  KFubKGj  )��}�(h�h�j  ]�j  KEj  KGubKHj  )��}�(h�h�j  ]�j  KEj  KHubKIj  )��}�(h�h�j  ]�j  KEj  KIubKJj  )��}�(h�h�j  ]�j  KEj  KJubKKj  )��}�(h�h�j  ]�j  KEj  KKubKLj  )��}�(h�h�j  ]�j  KEj  KLubKMj  )��}�(h�h�j  ]�j  KEj  KMubKNj  )��}�(h�h�j  ]�j  KEj  KNubKOj  )��}�(h�h�j  ]�j  KEj  KOubuKF}�(K j  )��}�(h�h�j  ]�j  KFj  K ubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubK	j  )��}�(h�h�j  ]�j  KFj  K	ubK
j  )��}�(h�h�j  ]�j  KFj  K
ubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubKj  )��}�(h�h�j  ]�j  KFj  KubK j  )��}�(h�h�j  ]�j  KFj  K ubK!j  )��}�(h�h�j  ]�j  KFj  K!ubK"j  )��}�(h�h�j  ]�j  KFj  K"ubK#j  )��}�(h�h�j  ]�j  KFj  K#ubK$j  )��}�(h�h�j  ]�j  KFj  K$ubK%j  )��}�(h�h�j  ]�j  KFj  K%ubK&j  )��}�(h�h�j  ]�j  KFj  K&ubK'j  )��}�(h�h�j  ]�j  KFj  K'ubK(j  )��}�(h�h�j  ]�j  KFj  K(ubK)j  )��}�(h�h�j  ]�j  KFj  K)ubK*j  )��}�(h�h�j  ]�j  KFj  K*ubK+j  )��}�(h�h�j  ]�j  KFj  K+ubK,j  )��}�(h�h�j  ]�j  KFj  K,ubK-j  )��}�(h�h�j  ]�j  KFj  K-ubK.j  )��}�(h�h�j  ]�j  KFj  K.ubK/j  )��}�(h�h�j  ]�j  KFj  K/ubK0j  )��}�(h�h�j  ]�j  KFj  K0ubK1j  )��}�(h�h�j  ]�j  KFj  K1ubK2j  )��}�(h�h�j  ]�j  KFj  K2ubK3j  )��}�(h�h�j  ]�j  KFj  K3ubK4j  )��}�(h�h�j  ]�j  KFj  K4ubK5j  )��}�(h�h�j  ]�j  KFj  K5ubK6j  )��}�(h�h�j  ]�j  KFj  K6ubK7j  )��}�(h�h�j  ]�j  KFj  K7ubK8j  )��}�(h�h�j  ]�j  KFj  K8ubK9j  )��}�(h�h�j  ]�j  KFj  K9ubK:j  )��}�(h�h�j  ]�j  KFj  K:ubK;j  )��}�(h�h�j  ]�j  KFj  K;ubK<j  )��}�(h�h�j  ]�j  KFj  K<ubK=j  )��}�(h�h�j  ]�j  KFj  K=ubK>j  )��}�(h�h�j  ]�j  KFj  K>ubK?j  )��}�(h�h�j  ]�j  KFj  K?ubK@j  )��}�(h�h�j  ]�j  KFj  K@ubKAj  )��}�(h�h�j  ]�j  KFj  KAubKBj  )��}�(h�h�j  ]�j  KFj  KBubKCj  )��}�(h�h�j  ]�j  KFj  KCubKDj  )��}�(h�h�j  ]�j  KFj  KDubKEj  )��}�(h�h�j  ]�j  KFj  KEubKFj  )��}�(h�h�j  ]�j  KFj  KFubKGj  )��}�(h�h�j  ]�j  KFj  KGubKHj  )��}�(h�h�j  ]�j  KFj  KHubKIj  )��}�(h�h�j  ]�j  KFj  KIubKJj  )��}�(h�h�j  ]�j  KFj  KJubKKj  )��}�(h�h�j  ]�j  KFj  KKubKLj  )��}�(h�h�j  ]�j  KFj  KLubKMj  )��}�(h�h�j  ]�j  KFj  KMubKNj  )��}�(h�h�j  ]�j  KFj  KNubKOj  )��}�(h�h�j  ]�j  KFj  KOubuKG}�(K j  )��}�(h�h�j  ]�j  KGj  K ubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubK	j  )��}�(h�h�j  ]�j  KGj  K	ubK
j  )��}�(h�h�j  ]�j  KGj  K
ubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubKj  )��}�(h�h�j  ]�j  KGj  KubK j  )��}�(h�h�j  ]�j  KGj  K ubK!j  )��}�(h�h�j  ]�j  KGj  K!ubK"j  )��}�(h�h�j  ]�j  KGj  K"ubK#j  )��}�(h�h�j  ]�j  KGj  K#ubK$j  )��}�(h�h�j  ]�j  KGj  K$ubK%j  )��}�(h�h�j  ]�j  KGj  K%ubK&j  )��}�(h�h�j  ]�j  KGj  K&ubK'j  )��}�(h�h�j  ]�j  KGj  K'ubK(j  )��}�(h�h�j  ]�j  KGj  K(ubK)j  )��}�(h�h�j  ]�j  KGj  K)ubK*j  )��}�(h�h�j  ]�j  KGj  K*ubK+j  )��}�(h�h�j  ]�j  KGj  K+ubK,j  )��}�(h�h�j  ]�j  KGj  K,ubK-j  )��}�(h�h�j  ]�j  KGj  K-ubK.j  )��}�(h�h�j  ]�j  KGj  K.ubK/j  )��}�(h�h�j  ]�j  KGj  K/ubK0j  )��}�(h�h�j  ]�j  KGj  K0ubK1j  )��}�(h�h�j  ]�j  KGj  K1ubK2j  )��}�(h�h�j  ]�j  �      KGj  K2ubK3j  )��}�(h�h�j  ]�j  KGj  K3ubK4j  )��}�(h�h�j  ]�j  KGj  K4ubK5j  )��}�(h�h�j  ]�j  KGj  K5ubK6j  )��}�(h�h�j  ]�j  KGj  K6ubK7j  )��}�(h�h�j  ]�j  KGj  K7ubK8j  )��}�(h�h�j  ]�j  KGj  K8ubK9j  )��}�(h�h�j  ]�j  KGj  K9ubK:j  )��}�(h�h�j  ]�j  KGj  K:ubK;j  )��}�(h�h�j  ]�j  KGj  K;ubK<j  )��}�(h�h�j  ]�j  KGj  K<ubK=j  )��}�(h�h�j  ]�j  KGj  K=ubK>j  )��}�(h�h�j  ]�j  KGj  K>ubK?j  )��}�(h�h�j  ]�j  KGj  K?ubK@j  )��}�(h�h�j  ]�j  KGj  K@ubKAj  )��}�(h�h�j  ]�j  KGj  KAubKBj  )��}�(h�h�j  ]�j  KGj  KBubKCj  )��}�(h�h�j  ]�j  KGj  KCubKDj  )��}�(h�h�j  ]�j  KGj  KDubKEj  )��}�(h�h�j  ]�j  KGj  KEubKFj  )��}�(h�h�j  ]�j  KGj  KFubKGj  )��}�(h�h�j  ]�j  KGj  KGubKHj  )��}�(h�h�j  ]�j  KGj  KHubKIj  )��}�(h�h�j  ]�j  KGj  KIubKJj  )��}�(h�h�j  ]�j  KGj  KJubKKj  )��}�(h�h�j  ]�j  KGj  KKubKLj  )��}�(h�h�j  ]�j  KGj  KLubKMj  )��}�(h�h�j  ]�j  KGj  KMubKNj  )��}�(h�h�j  ]�j  KGj  KNubKOj  )��}�(h�h�j  ]�j  KGj  KOubuKH}�(K j  )��}�(h�h�j  ]�j  KHj  K ubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubK	j  )��}�(h�h�j  ]�j  KHj  K	ubK
j  )��}�(h�h�j  ]�j  KHj  K
ubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubKj  )��}�(h�h�j  ]�j  KHj  KubK j  )��}�(h�h�j  ]�j  KHj  K ubK!j  )��}�(h�h�j  ]�j  KHj  K!ubK"j  )��}�(h�h�j  ]�j  KHj  K"ubK#j  )��}�(h�h�j  ]�j  KHj  K#ubK$j  )��}�(h�h�j  ]�j  KHj  K$ubK%j  )��}�(h�h�j  ]�j  KHj  K%ubK&j  )��}�(h�h�j  ]�j  KHj  K&ubK'j  )��}�(h�h�j  ]�j  KHj  K'ubK(j  )��}�(h�h�j  ]�j  KHj  K(ubK)j  )��}�(h�h�j  ]�j  KHj  K)ubK*j  )��}�(h�h�j  ]�j  KHj  K*ubK+j  )��}�(h�h�j  ]�j  KHj  K+ubK,j  )��}�(h�h�j  ]�j  KHj  K,ubK-j  )��}�(h�h�j  ]�j  KHj  K-ubK.j  )��}�(h�h�j  ]�j  KHj  K.ubK/j  )��}�(h�h�j  ]�j  KHj  K/ubK0j  )��}�(h�h�j  ]�j  KHj  K0ubK1j  )��}�(h�h�j  ]�j  KHj  K1ubK2j  )��}�(h�h�j  ]�j  KHj  K2ubK3j  )��}�(h�h�j  ]�j  KHj  K3ubK4j  )��}�(h�h�j  ]�j  KHj  K4ubK5j  )��}�(h�h�j  ]�j  KHj  K5ubK6j  )��}�(h�h�j  ]�j  KHj  K6ubK7j  )��}�(h�h�j  ]�j  KHj  K7ubK8j  )��}�(h�h�j  ]�j  KHj  K8ubK9j  )��}�(h�h�j  ]�j  KHj  K9ubK:j  )��}�(h�h�j  ]�j  KHj  K:ubK;j  )��}�(h�h�j  ]�j  KHj  K;ubK<j  )��}�(h�h�j  ]�j  KHj  K<ubK=j  )��}�(h�h�j  ]�j  KHj  K=ubK>j  )��}�(h�h�j  ]�j  KHj  K>ubK?j  )��}�(h�h�j  ]�j  KHj  K?ubK@j  )��}�(h�h�j  ]�j  KHj  K@ubKAj  )��}�(h�h�j  ]�j  KHj  KAubKBj  )��}�(h�h�j  ]�j  KHj  KBubKCj  )��}�(h�h�j  ]�j  KHj  KCubKDj  )��}�(h�h�j  ]�j  KHj  KDubKEj  )��}�(h�h�j  ]�j  KHj  KEubKFj  )��}�(h�h�j  ]�j  KHj  KFubKGj  )��}�(h�h�j  ]�j  KHj  KGubKHj  )��}�(h�h�j  ]�j  KHj  KHubKIj  )��}�(h�h�j  ]�j  KHj  KIubKJj  )��}�(h�h�j  ]�j  KHj  KJubKKj  )��}�(h�h�j  ]�j  KHj  KKubKLj  )��}�(h�h�j  ]�j  KHj  KLubKMj  )��}�(h�h�j  ]�j  KHj  KMubKNj  )��}�(h�h�j  ]�j  KHj  KNubKOj  )��}�(h�h�j  ]�j  KHj  KOubuKI}�(K j  )��}�(h�h�j  ]�j  KIj  K ubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubK	j  )��}�(h�h�j  ]�j  KIj  K	ubK
j  )��}�(h�h�j  ]�j  KIj  K
ubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubKj  )��}�(h�h�j  ]�j  KIj  KubK j  )��}�(h�h�j  ]�j  KIj  K ubK!j  )��}�(h�h�j  ]�j  KIj  K!ubK"j  )��}�(h�h�j  ]�j  KIj  K"ubK#j  )��}�(h�h�j  ]�j  KIj  K#ubK$j  )��}�(h�h�j  ]�j  KIj  K$ubK%j  )��}�(h�h�j  ]�j  KIj  K%ubK&j  )��}�(h�h�j  ]�j  KIj  K&ubK'j  )��}�(h�h�j  ]�j  KIj  K'ubK(j  )��}�(h�h�j  ]�j  KIj  K(ubK)j  )��}�(h�h�j  ]�j  KIj  K)ubK*j  )��}�(h�h�j  ]�j  KIj  K*ubK+j  )��}�(h�h�j  ]�j  KIj  K+ubK,j  )��}�(h�h�j  ]�j  KIj  K,ubK-j  )��}�(h�h�j  ]�j  KIj  K-ubK.j  )��}�(h�h�j  ]�j  KIj  K.ubK/j  )��}�(h�h�j  ]�j  KIj  K/ubK0j  )��}�(h�h�j  ]�j  KIj  K0ubK1j  )��}�(h�h�j  ]�j  KIj  K1ubK2j  )��}�(h�h�j  ]�j  KIj  K2ubK3j  )��}�(h�h�j  ]�j  KIj  K3ubK4j  )��}�(h�h�j  ]�j  KIj  K4ubK5j  )��}�(h�h�j  ]�j  KIj  K5ubK6j  )��}�(h�h�j  ]�j  KIj  K6ubK7j  )��}�(h�h�j  ]�j  KIj  K7ubK8j  )��}�(h�h�j  ]�j  KIj  K8ubK9j  )��}�(h�h�j  ]�j  KIj  K9ubK:j  )��}�(h�h�j  ]�j  KIj  K:ubK;j  )��}�(h�h�j  ]�j  KIj  K;ubK<j  )��}�(h�h�j  ]�j  KIj  K<ubK=j  )��}�(h�h�j  ]�j  KIj  K=ubK>j  )��}�(h�h�j  ]�j  KIj  K>ubK?j  )��}�(h�h�j  ]�j  KIj  K?ubK@j  )��}�(h�h�j  ]�j  KIj  K@ubKAj  )��}�(h�h�j  ]�j  KIj  KAubKBj  )��}�(h�h�j  ]�j  KIj  KBubKCj  )��}�(h�h�j  ]�j  KIj  KCubKDj  )��}�(h�h�j  ]�j  KIj  KDubKEj  )��}�(h�h�j  ]�j  KIj  KEubKFj  )��}�(h�h�j  ]�j  KIj  KFubKGj  )��}�(h�h�j  ]�j  KIj  KGubKHj  )��}�(h�h�j  ]�j  KIj  KHubKIj  )��}�(h�h�j  ]�j  KIj  KIubKJj  )��}�(h�h�j  ]�j  KIj  KJubKKj  )��}�(h�h�j  ]�j  KIj  KKubKLj  )��}�(h�h�j  ]�j  KIj  KLubKMj  )��}�(h�h�j  ]�j  KIj  KMubKNj  )��}�(h�h�j  ]�j  KIj  KNubKOj  )��}�(h�h�j  ]�j  KIj  KOubuKJ}�(K j  )��}�(h�h�j  ]�j  KJj  K ubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubK	j  )��}�(h�h�j  ]�j  KJj  K	ubK
j  )��}�(h�h�j  ]�j  KJj  K
ubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubKj  )��}�(h�h�j  ]�j  KJj  KubK j  )��}�(h�h�j  ]�j  KJj  K ubK!j  )��}�(h�h�j  ]�j  KJj  K!ubK"j  )��}�(h�h�j  ]�j  KJj  K"ubK#j  )��}�(h�h�j  ]�j  KJj  K#ubK$j  )��}�(h�h�j  ]�j  KJj  K$ubK%j  )��}�(h�h�j  ]�j  KJj  K%ubK&j  )��}�(h�h�j  ]�j  KJj  K&ubK'j  )��}�(h�h�j  ]�j  KJj  K'ubK(j  )��}�(h�h�j  ]�j  KJj  K(ubK)j  )��}�(h�h�j  ]�j  KJj  K)ubK*j  )��}�(h�h�j  ]�j  KJj  K*ubK+j  )��}�(h�h�j  ]�j  KJj  K+ubK,j  )��}�(h�h�j  ]�j  KJj  K,ubK-j  )��}�(h�h�j  ]�j  KJj  K-ubK.j  )��}�(h�h�j  ]�j  KJj  K.ubK/j  )��}�(h�h�j  ]�j  KJj  K/ubK0j  )��}�(h�h�j  ]�j  KJj  K0ubK1j  )��}�(h�h�j  ]�j  KJj  K1ubK2j  )��}�(h�h�j  ]�j  KJj  K2ubK3j  )��}�(h�h�j  ]�j  KJj  K3ubK4j  )��}�(h�h�j  ]�j  KJj  K4ubK5j  )��}�(h�h�j  ]�j  KJj  K5ubK6j  )��}�(h�h�j  ]�j  KJj  K6ubK7j  )��}�(h�h�j  ]�j  KJj  K7ubK8j  )��}�(h�h�j  ]�j  KJj  K8ubK9j  )��}�(h�h�j  ]�j  KJj  K9ubK:j  )��}�(h�h�j  ]�j  KJj  K:ubK;j  )��}�(h�h�j  ]�j  KJj  K;ubK<j  )��}�(h�h�j  ]�j  KJj  K<ubK=j  )��}�(h�h�j  ]�j  KJj  K=ubK>j  )��}�(h�h�j  ]�j  KJj  K>ubK?j  )��}�(h�h�j  ]�j  KJj  K?ubK@j  )��}�(h�h�j  ]�j  KJj  K@ubKAj  )��}�(h�h�j  ]�j  KJj  KAubKBj  )��}�(h�h�j  ]�j  KJj  KBubKCj  )��}�(h�h�j  ]�j  KJj  KCubKDj  )��}�(h�h�j  ]�j  KJj  KDubKEj  )��}�(h�h�j  ]�j  KJj  KEubKFj  )��}�(h�h�j  ]�j  KJj  KFubKGj  )��}�(h�h�j  ]�j  KJj  KGubKHj  )��}�(h�h�j  ]�j  KJj  KHubKIj  )��}�(h�h�j  ]�j  KJj  KIubKJj  )��}�(h�h�j  ]�j  KJj  KJubKKj  )��}�(h�h�j  ]�j  KJj  KKubKLj  )��}�(h�h�j  ]�j  KJj  KLubKMj  )��}�(h�h�j  ]�j  KJj  KMubKNj  )��}�(h�h�j  ]�j  KJj  KNubKOj  )��}�(h�h�j  ]�j  KJj  KOubuKK}�(K j  )��}�(h�h�j  ]�j  KKj  K ubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubK	j  )��}�(h�h�j  ]�j  KKj  K	ubK
j  )��}�(h�h�j  ]�j  KKj  K
ubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubKj  )��}�(h�h�j  ]�j  KKj  KubK j  )��}�(h�h�j  ]�j  KKj  K ubK!j  )��}�(h�h�j  ]�j  KKj  K!ubK"j  )��}�(h�h�j  ]�j  KKj  K"ubK#j  )��}�(h�h�j  ]�j  KKj  K#ubK$j  )��}�(h�h�j  ]�j  KKj  K$ubK%j  )��}�(h�h�j  ]�j  KKj  K%ubK&j  )��}�(h�h�j  ]�j  KKj  K&ubK'j  )��}�(h�h�j  ]�j  KKj  K'ubK(j  )��}�(h�h�j  ]�j  KKj  K(ubK)j  )��}�(h�h�j  ]�j  KKj  K)ubK*j  )��}�(h�h�j  ]�j  KKj  K*ubK+j  )��}�(h�h�j  ]�j  KKj  K+ubK,j  )��}�(h�h�j  ]�j  KKj  K,ubK-j  )��}�(h�h�j  ]�j  KKj  K-ubK.j  )��}�(h�h�j  ]�j  KKj  K.ubK/j  )��}�(h�h�j  ]�j  KKj  K/ubK0j  )��}�(h�h�j  ]�j  KKj  K0ubK1j  )��}�(h�h�j  ]�j  KKj  K1ubK2j  )��}�(h�h�j  ]�j  KKj  K2ubK3j  )��}�(h�h�j  ]�j  KKj  K3ubK4j  )��}�(h�h�j  ]�j  KKj  K4ubK5j  )��}�(h�h�j  ]�j  KKj  K5ubK6j  )��}�(h�h�j  ]�j  KKj  K6ubK7j  )��}�(h�h�j  ]�j  KKj  K7ubK8j  )��}�(h�h�j  ]�j  KKj  K8ubK9j  )��}�(h�h�j  ]�j  KKj  K9ubK:j  )��}�(h�h�j  ]�j  KKj  K:ubK;j  )��}�(h�h�j  ]�j  KKj  K;ubK<j  )��}�(h�h�j  ]�j  KKj  K<ubK=j  )��}�(h�h�j  ]�j  KKj  K=ubK>j  )��}�(h�h�j  ]�j  KKj  K>ubK?j  )��}�(h�h�j  ]�j  KKj  K?ubK@j  )��}�(h�h�j  ]�j  KKj  K@ubKAj  )��}�(h�h�j  ]�j  KKj  KAubKBj  )��}�(h�h�j  ]�j  KKj  KBubKCj  )��}�(h�h�j  ]�j  KKj  KCubKDj  )��}�(h�h�j  ]�j  KKj  KDubKEj  )��}�(h�h�j  ]�j  KKj  KEubKFj  )��}�(h�h�j  ]�j  KKj  KFubKGj  )��}�(h�h�j  ]�j  KKj  KGubKHj  )��}�(h�h�j  ]�j  KKj  KHubKIj  )��}�(h�h�j  ]�j  KKj  KIubKJj  )��}�(h�h�j  ]�j  KKj  KJubKKj  )��}�(h�h�j  ]�j  KKj  KKubKLj  )��}�(h�h�j  ]�j  KKj  KLubKMj  )��}�(h�h�j  ]�j  KKj  KMubKNj  )��}�(h�h�j  ]�j  KKj  KNubKOj  )��}�(h�h�j  ]�j  KKj  KOubuKL}�(K j  )��}�(h�h�j  ]�j  KLj  K ubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubK	j  )��}�(h�h�j  ]�j  KLj  K	ubK
j  )��}�(h�h�j  ]�j  KLj  K
ubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubKj  )��}�(h�h�j  ]�j  KLj  KubK j  )��}�(h�h�j  ]�j  KLj  K ubK!j  )��}�(h�h�j  ]�j  KLj  K!ubK"j  )��}�(h�h�j  ]�j  KLj  K"ubK#j  )��}�(h�h�j  ]�j  KLj  K#ubK$j  )��}�(h�h�j  ]�j  KLj  K$ubK%j  )��}�(h�h�j  ]�j  KLj  K%ubK&j  )��}�(h�h�j  ]�j  KLj  K&ubK'j  )��}�(h�h�j  ]�j  KLj  K'ubK(j  )��}�(h�h�j  ]�j  KLj  K(ubK)j  )��}�(h�h�j  ]�j  KLj  K)ubK*j  )��}�(h�h�j  ]�j  KLj  K*ubK+j  )��}�(h�h�j  ]�j  KLj  K+ubK,j  )��}�(h�h�j  ]�j  KLj  K,ubK-j  )��}�(h�h�j  ]�j  KLj  K-ubK.j  )��}�(h�h�j  ]�j  KLj  K.ubK/j  )��}�(h�h�j  ]�j  KLj  K/ubK0j  )��}�(h�h�j  ]�j  KLj  K0ubK1j  )��}�(h�h�j  ]�j  KLj  K1ubK2j  )��}�(h�h�j  ]�j  KLj  K2ubK3j  )��}�(h�h�j  ]�j  KLj  K3ubK4j  )��}�(h�h�j  ]�j  KLj  K4ubK5j  )��}�(h�h�j  ]�j  KLj  K5ubK6j  )��}�(h�h�j  ]�j  KLj  K6ubK7j  )��}�(h�h�j  ]�j  KLj  K7ubK8j  )��}�(h�h�j  ]�j  KLj  K8ubK9j  )��}�(h�h�j  ]�j  KLj  K9ubK:j  )��}�(h�h�j  ]�j  KLj  K:ubK;j  )��}�(h�h�j  ]�j  KLj  K;ubK<j  )��}�(h�h�j  ]�j  KLj  K<ubK=j  )��}�(h�h�j  ]�j  KLj  K=ubK>j  )��}�(h�h�j  ]�j  KLj  K>ubK?j  )��}�(h�h�j  ]�j  KLj  K?ubK@j  )��}�(h�h�j  ]�j  KLj  K@ubKAj  )��}�(h�h�j  ]�j  KLj  KAubKBj  )��}�(h�h�j  ]�j  KLj  KBubKCj  )��}�(h�h�j  ]�j  KLj  KCubKDj  )��}�(h�h�j  ]�j  KLj  KDubKEj  )��}�(h�h�j  ]�j  KLj  KEubKFj  )��}�(h�h�j  ]�j  KLj  KFubKGj  )��}�(h�h�j  ]�j  KLj  KGubKHj  )��}�(h�h�j  ]�j  KLj  KHubKIj  )��}�(h�h�j  ]�j  KLj  KIubKJj  )��}�(h�h�j  ]�j  KLj  KJubKKj  )��}�(h�h�j  ]�j  KLj  KKubKLj  )��}�(h�h�j  ]�j  KLj  KLubKMj  )��}�(h�h�j  ]�j  KLj  KMubKNj  )��}�(h�h�j  ]�j  KLj  KNubKOj  )��}�(h�h�j  ]�j  KLj  KOubuKM}�(K j  )��}�(h�h�j  ]�j  KMj  K ubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubK	j  )��}�(h�h�j  ]�j  KMj  K	ubK
j  )��}�(h�h�j  ]�j  KMj  K
ubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubKj  )��}�(h�h�j  ]�j  KMj  KubK j  )��}�(h�h�j  ]�j  KMj  K ubK!j  )��}�(h�h�j  ]�j  KMj  K!ubK"j  )��}�(h�h�j  ]�j  KMj  K"ubK#j  )��}�(h�h�j  ]�j  KMj  K#ubK$j  )��}�(h�h�j  ]�j  KMj  K$ubK%j  )��}�(h�h�j  ]�j  KMj  K%ubK&j  )��}�(h�h�j  ]�j  KMj  K&ubK'j  )��}�(h�h�j  ]�j  KMj  K'ubK(j  )��}�(h�h�j  ]�j  KMj  K(ubK)j  )��}�(h�h�j  ]�j  KMj  K)ubK*j  )��}�(h�h�j  ]�j  KMj  K*ubK+j  )��}�(h�h�j  ]�j  KMj  K+ubK,j  )��}�(h�h�j  ]�j  KMj  K,ubK-j  )��}�(h�h�j  ]�j  KMj  K-ubK.j  )��}�(h�h�j  ]�j  KMj  K.ubK/j  )��}�(h�h�j  ]�j  KMj  K/ubK0j  )��}�(h�h�j  ]�j  KMj  K0ubK1j  )��}�(h�h�j  ]�j  KMj  K1ubK2j  )��}�(h�h�j  ]�j  KMj  K2ubK3j  )��}�(h�h�j  ]�j  KMj  K3ubK4j  )��}�(h�h�j  ]�j  KMj  K4ubK5j  )��}�(h�h�j  ]�j  KMj  K5ubK6j  )��}�(h�h�j  ]�j  KMj  K6ubK7j  )��}�(h�h�j  ]�j  KMj  K7ubK8j  )��}�(h�h�j  ]�j  KMj  K8ubK9j  )��}�(h�h�j  ]�j  KMj  K9ubK:j  )��}�(h�h�j  ]�j  KMj  K:ubK;j  )��}�(h�h�j  ]�j  KMj  K;ubK<j  )��}�(h�h�j  ]�j  KMj  K<ubK=j  )��}�(h�h�j  ]�j  KMj  K=ubK>j  )��}�(h�h�j  ]�j  KMj  K>ubK?j  )��}�(h�h�j  ]�j  KMj  K?ubK@j  )��}�(h�h�j  ]�j  KMj  K@ubKAj  )��}�(h�h�j  ]�j  KMj  KAubKBj  )��}�(h�h�j  ]�j  KMj  KBubKCj  )��}�(h�h�j  ]�j  KMj  KCubKDj  )��}�(h�h�j  ]�j  KMj  KDubKEj  )��}�(h�h�j  ]�j  KMj  KEubKFj  )��}�(h�h�j  ]�j  KMj  KFubKGj  )��}�(h�h�j  ]�j  KMj  KGubKHj  )��}�(h�h�j  ]�j  KMj  KHubKIj  )��}�(h�h�j  ]�j  KMj  KIubKJj  )��}�(h�h�j  ]�j  KMj  KJubKKj  )��}�(h�h�j  ]�j  KMj  KKubKLj  )��}�(h�h�j  ]�j  KMj  KLubKMj  )��}�(h�h�j  ]�j  KMj  KMubKNj  )��}�(h�h�j  ]�j  KMj  KNubKOj  )��}�(h�h�j  ]�j  KMj  KOubuKN}�(K j  )��}�(h�h�j  ]�j  KNj  K ubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubK	j  )��}�(h�h�j  ]�j  KNj  K	ubK
j  )��}�(h�h�j  ]�j  KNj  K
ubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubKj  )��}�(h�h�j  ]�j  KNj  KubK j  )��}�(h�h�j  ]�j  KNj  K ubK!j  )��}�(h�h�j  ]�j  KNj  K!ubK"j  )��}�(h�h�j  ]�j  KNj  K"ubK#j  )��}�(h�h�j  ]�j  KNj  K#ubK$j  )��}�(h�h�j  ]�j  KNj  K$ubK%j  )��}�(h�h�j  ]�j  KNj  K%ubK&j  )��}�(h�h�j  ]�j  KNj  K&ubK'j  )��}�(h�h�j  ]�j  KNj  K'ubK(j  )��}�(h�h�j  ]�j  KNj  K(ubK)j  )��}�(h�h�j  ]�j  KNj  K)ubK*j  )��}�(h�h�j  ]�j  KNj  K*ubK+j  )��}�(h�h�j  ]�j  KNj  K+ubK,j  )��}�(h�h�j  ]�j  KNj  K,ubK-j  )��}�(h�h�j  ]�j  KNj  K-ubK.j  )��}�(h�h�j  ]�j  KNj  K.ubK/j  )��}�(h�h�j  ]�j  KNj  K/ubK0j  )��}�(h�h�j  ]�j  KNj  K0ubK1j  )��}�(h�h�j  ]�j  KNj  K1ubK2j  )��}�(h�h�j  ]�j  KNj  K2ubK3j  )��}�(h�h�j  ]�j  KNj  K3ubK4j  )��}�(h�h�j  ]�j  KNj  K4ubK5j  )��}�(h�h�j  ]�j  KNj  K5ubK6j  )��}�(h�h�j  ]�j  KNj  K6ubK7j  )��}�(h�h�j  ]�j  KNj  K7ubK8j  )��}�(h�h�j  ]�j  KNj  K8ubK9j  )��}�(h�h�j  ]�j  KNj  K9ubK:j  )��}�(h�h�j  ]�j  KNj  K:ubK;j  )��}�(h�h�j  ]�j  KNj  K;ubK<j  )��}�(h�h�j  ]�j  KNj  K<ubK=j  )��}�(h�h�j  ]�j  KNj  K=ubK>j  )��}�(h�h�j  ]�j  KNj  K>ubK?j  )��}�(h�h�j  ]�j  KNj  K?ubK@j  )��}�(h�h�j  ]�j  KNj  K@ubKAj  )��}�(h�h�j  ]�j  KNj  KAubKBj  )��}�(h�h�j  ]�j  KNj  KBubKCj  )��}�(h�h�j  ]�j  KNj  KCubKDj  )��}�(h�h�j  ]�j  KNj  KDubKEj  )��}�(h�h�j  ]�j  KNj  KEubKFj  )��}�(h�h�j  ]�j  KNj  KFubKGj  )��}�(h�h�j  ]�j  KNj  KGubKHj  )��}�(h�h�j  ]�j  KNj  KHubKIj  )��}�(h�h�j  ]�j  KNj  KIubKJj  )��}�(h�h�j  ]�j  KNj  KJubKKj  )��}�(h�h�j  ]�j  KNj  KKubKLj  )��}�(h�h�j  ]�j  KNj  KLubKMj  )��}�(h�h�j  ]�j  KNj  KMubKNj  )��}�(h�h�j  ]�j  KNj  KNubKOj  )��}�(h�h�j  ]�j  KNj  KOubuKO}�(K j  )��}�(h�h�j  ]�j  KOj  K ubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubK	j  )��}�(h�h�j  ]�j  KOj  K	ubK
j  )��}�(h�h�j  ]�j  KOj  K
ubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubKj  )��}�(h�h�j  ]�j  KOj  KubK j  )��}�(h�h�j  ]�j  KOj  K ubK!j  )��}�(h�h�j  ]�j  KOj  K!ubK"j  )��}�(h�h�j  ]�j  KOj  K"ubK#j  )��}�(h�h�j  ]�j  KOj  K#ubK$j  )��}�(h�h�j  ]�j  KOj  K$ubK%j  )��}�(h�h�j  ]�j  KOj  K%ubK&j  )��}�(h�h�j  ]�j  KOj  K&ubK'j  )��}�(h�h�j  ]�j  KOj  K'ubK(j  )��}�(h�h�j  ]�j  KOj  K(ubK)j  )��}�(h�h�j  ]�j  KOj  K)ubK*j  )��}�(h�h�j  ]�j  KOj  K*ubK+j  )��}�(h�h�j  ]�j  KOj  K+ubK,j  )��}�(h�h�j  ]�j  KOj  K,ubK-j  )��}�(h�h�j  ]�j  KOj  K-ubK.j  )��}�(h�h�j  ]�j  KOj  K.ubK/j  )��}�(h�h�j  ]�j  KOj  K/ubK0j  )��}�(h�h�j  ]�j  KOj  K0ubK1j  )��}�(h�h�j  ]�j  KOj  K1ubK2j  )��}�(h�h�j  ]�j  KOj  K2ubK3j  )��}�(h�h�j  ]�j  KOj  K3ubK4j  )��}�(h�h�j  ]�j  KOj  K4ubK5j  )��}�(h�h�j  ]�j  KOj  K5ubK6j  )��}�(h�h�j  ]�j  KOj  K6ubK7j  )��}�(h�h�j  ]�j  KOj  K7ubK8j  )��}�(h�h�j  ]�j  KOj  K8ubK9j  )��}�(h�h�j  ]�j  KOj  K9ubK:j  )��}�(h�h�j  ]�j  KOj  K:ubK;j  )��}�(h�h�j  ]�j  KOj  K;ubK<j  )��}�(h�h�j  ]�j  KOj  K<ubK=j  )��}�(h�h�j  ]�j  KOj  K=ubK>j  )��}�(h�h�j  ]�j  KOj  K>ubK?j  )��}�(h�h�j  ]�j  KOj  K?ubK@j  )��}�(h�h�j  ]�j  KOj  K@ubKAj  )��}�(h�h�j  ]�j  KOj  KAubKBj  )��}�(h�h�j  ]�j  KOj  KBubKCj  )��}�(h�h�j  ]�j  KOj  KCubKDj  )��}�(h�h�j  ]�j  KOj  KDubKEj  )��}�(h�h�j  ]�j  KOj  KEubKFj  )��}�(h�h�j  ]�j  KOj  KFubKGj  )��}�(h�h�j  ]�j  KOj  KGubKHj  )��}�(h�h�j  ]�j  KOj  KHubKIj  )��}�(h�h�j  ]�j  KOj  KIubKJj  )��}�(h�h�j  ]�j  KOj  KJubKKj  )��}�(h�h�j  ]�j  KOj  KKubKLj  )��}�(h�h�j  ]�j  KOj  KLubKMj  )��}�(h�h�j  ]�j  KOj  KMubKNj  )��}�(h�h�j  ]�j  KOj  KNubKOj  )��}�(h�h�j  ]�j  KOj  KOubuu�	enemyList�]�(j  j�  e�master_Changed_Tiles�]�(]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KEKe]�(KDKe]�(KEKe]�(KDKe]�(KEKe]�(KDKe]�(KEKe]�(KDKe]�(KEKe]�(KDKe]�(KEKe]�(KDKe]�(KEKe]�(KEKe]�(KDKe]�(KEKe]�(KEKe]�(KDKe]�(KEKe]�(KEKe]�(KEKe]�(KDKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KDKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KDKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEK
e]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KFKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KFKe]�(KEKe]�(KEKe]�(KFKe]�(KEKe]�(KEKe]�(KEKe]�(KFKe]�(KEKe]�(KFKe]�(KEKe]�(KEKe]�(KFKe]�(KEKe]�(KFKe]�(KEKe]�(KFKe]�(KEKe]�(KFKe]�(KEKe]�(KFKe]�(KFKe]�(KEKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKeeh[hԌdjikstra_Player�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�P�     G�P�     G�P      G�P�     G�P�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�P�     G�P      G�O�     G�P      G�P�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�P      G�O�     G�N�     G�O�     G�P      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�O�     G�N�     G�N      G�N�     G�O�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�N�     G�N      G�M@     G�N      G�N�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�N      G�M@     G�L�     G�M@     G�N      G�N�     G�O�     G�P      G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      G�S�     G�S�     G�T@     NNNNNNNNNNNNG�U`     G�U      G�T�     G�T@     G�S�     G�T@     G�T�     G�U      G�U`     G�U�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�M@     G�L�     G�K�     G�L�     G�M@     NNNNNNNNNNNNNG�T�     NNNNNNNNNNNNG�U      G�T�     G�T@     G�S�     G�S�     G�S�     G�T@     G�T�     G�U      G�U`     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�L�     G�K�     G�K      G�K�     G�L�     NNNNNNNNNNNNNG�U      NNNNNNNNNNNNNNNNG�S      G�S�     G�S�     G�T@     G�T�     G�U      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�J@     G�K      G�K�     NNNNNNNNNNNNNG�U`     NNNNNNNNNNNNNNNNG�R�     G�S      G�S�     G�S�     G�T@     G�T�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�I�     G�J@     G�K      NNNNNNNNNNNNNG�U�     NNNNNNNNNNNNNNNNG�R`     G�R�     G�S      G�S�     G�S�     G�T@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�H�     NNNNNNNNNNNNNNNG�V      NNNNNNNNNNNNNG�Q�     NNG�R      G�R`     G�R�     G�S      G�S�     G�S�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�H      NNNNNNNNNNNNNNNK NNNNNNNNNNNNG�Q�     G�Q@     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      G�S�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�G@     NNNNNNNNNNNNNNNG�V      NNNNNNNNNNNNG�Q@     G�P�     G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�F�     NNNNNNNNNNNNNNNG�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�E�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�O�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�B�     G�C�     G�D@     G�E      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�N�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�B      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�N      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�A@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�M@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�@�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�L�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�?�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�K�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�>      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�K      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�<�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�J@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�;      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�I�     G�J@     G�K      G�K�     G�L�     G�M@     G�N      G�N�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�>      G�<�     G�;      G�9�     G�8      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�H�     G�I�     G�J@     G�K      G�K�     G�L�     G�M@     G�N      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�<�     G�;      G�9�     G�8      G�6�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�H      G�H�     G�I�     G�J@     G�K      G�K�     G�L�     G�M@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�;      G�9�     G�8      G�6�     G�5      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�G@     G�H      G�H�     G�I�     G�J@     G�K      G�K�     G�L�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�9�     G�8      G�6�     G�5      G�3�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�F�     G�G@     G�H      G�H�     G�I�     G�J@     G�K      G�K�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�8      G�6�     G�5      G�3�     G�2      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�E�     G�F�     G�G@     G�H      G�H�     G�I�     G�J@     G�K      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�6�     G�5      G�3�     G�2      G�0�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�E      G�E�     G�F�     G�G@     G�H      G�H�     G�I�     G�J@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�5      G�3�     G�2      G�0�     G�.      NNNNNNNNNNNNNNNG�.      G�0�     G�2      G�3�     G�5      G�6�     G�8      G�9�     G�;      G�<�     G�>      G�?�     G�@�     G�A@     G�B      G�B�     G�C�     G�D@     G�E      G�E�     G�F�     G�G@     G�H      G�H�     G�I�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNG�0�     G�.      G�+      NNNNNNNNNNNNNNNG�+      NNNNNNNNNNNNNNNNNG�E�     G�F�     G�G@     G�H      G�H�     G�I�     G�J@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNG�.      G�+      G�(      G�%      G�"      G�      G�      G�      G�      G��      G�       G��      G�      G�      G�      G�      G�"      G�%      G�(      NNNNNNNNNNNNNNNNNNG�G@     G�H      G�H�     G�I�     G�J@     G�K      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�	decorList�]�(j�  jo  j  e�	textSpace��Ornate mosaic floor
��SeenMap�]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K ee�maze�]�(]�(�#�j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  �.�j�O  j~  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  jl  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jl  jl  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jl  jl  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  hUj�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jl  jl  j�O  j�O  j�O  j�  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  �      j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jA  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jl  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jM  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jM  jM  jM  jM  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jM  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  hUj�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  h0j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jM  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jM  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jl  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  ee�levelManager��LevelManager�jP  ��)��}�(�nextSeed�M&�	levelList�]�(h�)��}�(h�Kh�]�(KKKKKKeh�]�(hQh�h�h�hrh�h�h�hbhlh�h�h�h�h<h�h�h%h�h]h�h�eh�]�hQah�]�(h�h�h�hbhlh�h�h�h�h<h�h�h%h�h]h�h�eh�]�(KKeh�h�j  }�(K h�)��}�(h�jP  h/jl  j  K j  Kj  Kh�j�  )��}�(h2j�  h[jP  h/jl  ubh2j�  ubKh�)��}�(h�jP  h/jM  j  Kj  Kj  Kh�jO  )��}�(h[jP  h-jR  h/jM  h2jN  ubh2jN  ubKh�)��}�(h�jP  h/hUj  Kj  Kj  K"h�hQ)��}�(h)�h*�hTKh[jP  h,h*h-h.h/hUh2hVubh2j  ubKh�)��}�(h�jP  h/jM  j  Kj  Kj  Kh�jO  )��}�(h[j!P  h-jR  h/jM  h2jN  ubh2jN  ubKh�)��}�(h�jP  h/jM  j  Kj  Kj  Kh�jP  )��}�(hM]�(h�)��}�(�
arrowCount�Kh*�h,h*h-h.h/�i�h)�h2�Bundle of Arrows�ubh�)��}�(hKh)�h*�huhh,hvh-h.h/hwh2�Scroll of Fireball�ubh�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2�Leather Shirt�ubjb  )��}�(h)�h*�h,h*h-je  h/jf  jg  K	h2jh  ubeh[j%P  h-ji  h/jM  h2jO  ubh2jO  ubKh�)��}�(h�jP  h/j  j  Kj  Kj  K h�j�  )��}�(hKhK h/j  j  K(j  ]�(j7P  h�)��}�(h�jP  h/j  j  K	j  Kj  K%h�j  )��}�(hKhK h/j  j  K(j  ]�(j7P  j<P  eh Kh!�h"h%)��}�(h(K
hKh)�h*�h+Kh,h"h-h.h/h0h1�h2h3ubh4K h5Kh6K h7K h8K	h9Kh�Kh@Nj#  G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2j4P  ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4Kh1�h2hkubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j<P  j/  Kdj0  ]�j2  K h-j3  h2j  ubh2j4  ubeh Kh!�h"h])��}�(h(KhKh)�h*�h+Kh,h"h-h.h/h0h1�h2h`ubh4K h5Kh6K h7K h8Kh9Kh�Kh@hb)��}�(hKh/h0h,heh)�h*�hG�h(Kh K h+KhIK h-h.hHKhJ�h1�h2hfubj#  G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2j4P  ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4Kh1�h2hkubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j7P  j/  Kdj0  ]�j2  K h-j3  h2j�  ubh2j4  ubKh�)��}�(h�jP  h/jA  j  Kj  Kj  Kh�jC  )��}�(h[jUP  h�jP  j�  Kj  J����j  Kj  Kh�Nh2j�  ubh2jF  ubKh�)��}�(h�jP  h/h�j  Kj  K(j  K)h�hh2h ubKh�)��}�(h�jP  h/jl  j  Kj  Kj  Kh�j  )��}�(h2j  h[j[P  h/jl  ubh2j  ubK	j<P  K
h�)��}�(h�jP  h/j  j  K
j  Kj  Kh�j  )��}�(hKhK h/j  j  K(j  ]�(j_P  h�)��}�(h�jP  h/j  j  Kj  Kj  K"h�j  )��}�(hKhK h/j  j  K(j  ]�(j_P  jdP  eh Kh!�h"h%)��}�(h(K
hKh)�h*�h+Kh,h"h-h.h/h0h1�h2h3ubh4K h5Kh6K h7K h8K	h9Kh�Kh@Nj#  G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2j4P  ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4Kh1�h2hkubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[jdP  j/  Kdj0  ]�j2  K h-j3  h2j  ubh2j4  ubeh Kh!�h"h%)��}�(h(K
hKh)�h*�h+Kh,h"h-h.h/h0h1�h2h3ubh4K h5Kh6K h7K h8K	h9Kh�Kh@Nj#  G        hK�hL�hM]�h:h�)��}�(h(KhKh)�h*�h+Kh,h:h-h.h/h0h1�h2j4P  ubhHKh��h�Nh�K h�Nh�hl)��}�(hKh/h0h,heh)�h*�hG�hHKh Kh+KhIKhJ�h-h.h4Kh1�h2hkubj*  Nh(K j+  �hh�K j,  Nh�Kj-  Kh�Nh͉h�]�h[j_P  j/  Kdj0  ]�j2  K h-j3  h2j  ubh2j4  ubKjdP  Kh�)��}�(h�jP  h/jM  j  Kj  Kj  K	h�jP  )��}�(hM]�h[j{P  h-h.h/jM  h2jO  ubh2jO  ubKh�)��}�(h�jP  h/hUj  Kj  K!j  Kh�hyh2j  ubKh�)��}�(h�jP  h/jl  j  Kj  K(j  K%h�j�  )��}�(h2j�  h[j�P  h/jl  ubh2j�  ubKh�)��}�(h�jP  h/j~  j  Kj  K(j  K)h�j�  )��}�(h�jP  h[j�P  j  J����j  K(j�  Kh�Nj  K)h2j�  ubh2j�  ubKh�)��}�(h�jP  h/jM  j  Kj  K)j  K'h�jP  )��}�(hM]�h[j�P  h-h.h/jM  h2jO  ubh2jO  ubKh�)��}�(h�jP  h/jM  j  Kj  K-j  K%h�jP  )��}�(hM]�h[j�P  h-h.h/jM  h2jO  ubh2jO  ubKh�)��}�(h�jP  h/h0j  Kj  Kj  K	h�hYh2h3ubKh�)��}�(h�jP  h/h0j  Kj  Kj  K	h�hoh2hkubKh�)��}�(h�jP  h/h0j  Kj  Kj  Kh�hih2h`ubKh�)��}�(h�jP  h/h0j  Kj  Kj  Kh�hmh2hkubKh�)��}�(h�jP  h/hwj  Kj  Kj  Kh�hsh2hxubKh�)��}�(h�jP  h/h0j  Kj  K*j  Kh�h{h2h`ubKh�)��}�(h�jP  h/h0j  Kj  K*j  Kh�h}h2hkubKh�)��}�(h�jP  h/jf  j  Kj  K*j  Kh�jb  )��}�(h)�h*�h[Nh,h*h-je  h/jf  jg  Kh2jh  ubh2jh  ubKh�)��}�(h�jP  h/h0j  Kj  K,j  K$h�hh2h`ubK h�)��}�(h�jP  h/h0j  K j  K,j  K$h�h�h2hkubK!h�)��}�(h�jP  h/jf  j  K!j  K,j  K$h�jb  )��}�(h)�h*�h[Nh,h*h-je  h/jf  jg  Kh2jh  ubh2jh  ubK"h�)��}�(h�jP  h/h0j  K"j  K+j  K$h�h�h2h`ubK#h�)��}�(h�jP  h/h0j  K#j  K+j  K$h�h�h2hkubK$h�)��}�(h�jP  h/h�j  K$j  K+j  K$h�h�h2h�ubujk  ]�(]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKK K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKKK K K K K KKKKKKKKKKKK KKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKKKKKKKKKK KKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKKKKKKKKKK KKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKKKKKKKKKK KKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKK K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKK KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKK KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKK KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKK KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K K K K K K K K K K K KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKK K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKeej�  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNK[KZKYKZNNNNNNNNNNNKfKgKhKiKjKkKlKmKnKoKpKqKpKoKnKoKpKqKrNNNNNNNNNNNNNNNNNNNNNNe]�(NNNK[KZKYKXKYNNNNNNNNNNNKeNNNNNNNNNNKpKoKnKmKnKoKpKqNNNNNNNNNNNNNNNNNNNNNNe]�(NNK[KZKYKXKWKXNNNNNNNNNNNKdNNNNNNNNNNKoKnKmKlKmKnKoKpNNNNNNNNNNNNNNNNNNNNNNe]�(NNKZKYKXKWKVKWNNNNNNNNNNNKcNNNNNNNNNNKnKmKlKkKlKmKnKoNNNNNNNNNNNNNNNNNNNNNNe]�(NNKYKXKWKVKUKVNNNNNNNNNNNKbNNNNNNNNNNNKlKkKjKkKlKmKnNNNNNNNNNNNNNNNNNNNNNNe]�(NNKXKWKVKUKTKUKVKWKXKYKZK[K\K]K^K_K`KaNNNNNNNNNNNNKjKiKjKkKlKmNNNNNNNNNNNNNNNNNNNNNNe]�(NNKWKVKUKTKSKTNNNNNNNNNNNNNNNNNNNNNNNNNKhNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKVKUKTKSKRKSNNNNNNNNNNNNNNNNNNNNNNNNNKgNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKUKTKSKRKQKRNNNNNNNNNNNNNNNNNNNNNNNNNKfNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKPNNNNNNNNNNNNNNNNNNNNNNNNNNKeNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKONNNNNNNNNNNNNNNNNNNNNNNNNNKdNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNKcNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKMNNNNNNNNNNNNNNNNNNNNNNNNNNKbNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKLNNNNNNNNNNNNNNNNNNNNNNNNNNKaNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKKKJKIKHNNNNNNNNNNNNNNNNNNNNNNNK`NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNNNNK_NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNNNNK^NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKENNNNNNNNNNNNNNNNNNNNNNNK]NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNNNNK\NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNNNNK[NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKBNNNNNNNNNNNNNKPKQKRKSKTKUKVKWKXKYKZK[K\K]NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKANNNNNNNNNNNNNKONNNNNNKXKYKZK[K\K]K^NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK>K?K@KAKBKCNNNNNNNNNNKNNNNNNNKYKZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK=K>K?K@KAKBNNNNNNNNNNKMNNNNNNKZK[K\K]K^K_K`NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK<K=K>K?K@KANNNNNNNNNNKLNNNNNNK[K\K]K^K_K`KaNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK;K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKNNNNNNK\K]K^K_K`KaKbNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK:K;K<K=K>K?NNNNNNNNNNNNNNNNNK]K^K_K`KaKbKcNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK9K:K;K<K=K>NNNNNNNNNNNNNNNNNK^K_K`KaKbKcKdNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK8K9K:K;K<K=NNNNNNNNNNNNNNNNNK_K`KaKbKcKdKeNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK7K8K9K:K;K<NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK6NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK5NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK4NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK3NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNK.K/K0K1NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK-NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKK NNNNNNNNNNNNNNNNNNe]�(NNNNK,NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK+K*K)K(K'NNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK*K)K(K'K&K%K$K#K"K!K KKKKKNNNNNNNNNNNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK+K*K)K(K'NNNNNNNNNNKKKKKKKKKKKKKKKKK
K	KKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK,K+K*K)K(NNNNNNNNNNNNNNNNNNNNNNNNNNNK
K	KKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK-K,K+K*K)NNNNNNNNNNNNNNNNNNNNNNNNNNNKK
K	KKKNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKK
K	KKNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej  }�(K }�(K j  )��}�(h�jP  j  ]�j  K j  K ubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubK	j  )��}�(h�jP  j  ]�j  K j  K	ubK
j  )��}�(h�jP  j  ]�j  K j  K
ubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubK j  )��}�(h�jP  j  ]�j  K j  K ubK!j  )��}�(h�jP  j  ]�j  K j  K!ubK"j  )��}�(h�jP  j  ]�j  K j  K"ubK#j  )��}�(h�jP  j  ]�j  K j  K#ubK$j  )��}�(h�jP  j  ]�j  K j  K$ubK%j  )��}�(h�jP  j  ]�j  K j  K%ubK&j  )��}�(h�jP  j  ]�j  K j  K&ubK'j  )��}�(h�jP  j  ]�j  K j  K'ubK(j  )��}�(h�jP  j  ]�j  K j  K(ubK)j  )��}�(h�jP  j  ]�j  K j  K)ubK*j  )��}�(h�jP  j  ]�j  K j  K*ubK+j  )��}�(h�jP  j  ]�j  K j  K+ubK,j  )��}�(h�jP  j  ]�j  K j  K,ubK-j  )��}�(h�jP  j  ]�j  K j  K-ubK.j  )��}�(h�jP  j  ]�j  K j  K.ubK/j  )��}�(h�jP  j  ]�j  K j  K/ubK0j  )��}�(h�jP  j  ]�j  K j  K0ubK1j  )��}�(h�jP  j  ]�j  K j  K1ubK2j  )��}�(h�jP  j  ]�j  K j  K2ubK3j  )��}�(h�jP  j  ]�j  K j  K3ubK4j  )��}�(h�jP  j  ]�j  K j  K4ubK5j  )��}�(h�jP  j  ]�j  K j  K5ubK6j  )��}�(h�jP  j  ]�j  K j  K6ubK7j  )��}�(h�jP  j  ]�j  K j  K7ubK8j  )��}�(h�jP  j  ]�j  K j  K8ubK9j  )��}�(h�jP  j  ]�j  K j  K9ubK:j  )��}�(h�jP  j  ]�j  K j  K:ubK;j  )��}�(h�jP  j  ]�j  K j  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�K aj  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�Kaj  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�Kaj  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�Kaj  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�Kaj  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�Kaj  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�Kaj  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�Kaj  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�K	aj  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK	}�(K j  )��}�(h�jP  j  ]�j  K	j  K ubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubK	j  )��}�(h�jP  j  ]�j  K	j  K	ubK
j  )��}�(h�jP  j  ]�j  K	j  K
ubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubKj  )��}�(h�jP  j  ]�j  K	j  KubK j  )��}�(h�jP  j  ]�j  K	j  K ubK!j  )��}�(h�jP  j  ]�j  K	j  K!ubK"j  )��}�(h�jP  j  ]�j  K	j  K"ubK#j  )��}�(h�jP  j  ]�j  K	j  K#ubK$j  )��}�(h�jP  j  ]�j  K	j  K$ubK%j  )��}�(h�jP  j  ]�j  K	j  K%ubK&j  )��}�(h�jP  j  ]�j  K	j  K&ubK'j  )��}�(h�jP  j  ]�j  K	j  K'ubK(j  )��}�(h�jP  j  ]�j  K	j  K(ubK)j  )��}�(h�jP  j  ]�j  K	j  K)ubK*j  )��}�(h�jP  j  ]�j  K	j  K*ubK+j  )��}�(h�jP  j  ]�j  K	j  K+ubK,j  )��}�(h�jP  j  ]�j  K	j  K,ubK-j  )��}�(h�jP  j  ]�j  K	j  K-ubK.j  )��}�(h�jP  j  ]�j  K	j  K.ubK/j  )��}�(h�jP  j  ]�j  K	j  K/ubK0j  )��}�(h�jP  j  ]�j  K	j  K0ubK1j  )��}�(h�jP  j  ]�j  K	j  K1ubK2j  )��}�(h�jP  j  ]�j  K	j  K2ubK3j  )��}�(h�jP  j  ]�j  K	j  K3ubK4j  )��}�(h�jP  j  ]�j  K	j  K4ubK5j  )��}�(h�jP  j  ]�j  K	j  K5ubK6j  )��}�(h�jP  j  ]�j  K	j  K6ubK7j  )��}�(h�jP  j  ]�j  K	j  K7ubK8j  )��}�(h�jP  j  ]�j  K	j  K8ubK9j  )��}�(h�jP  j  ]�j  K	j  K9ubK:j  )��}�(h�jP  j  ]�j  K	j  K:ubK;j  )��}�(h�jP  j  ]�j  K	j  K;ubuK
}�(K j  )��}�(h�jP  j  ]�j  K
j  K ubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubK	j  )��}�(h�jP  j  ]�j  K
j  K	ubK
j  )��}�(h�jP  j  ]�j  K
j  K
ubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubKj  )��}�(h�jP  j  ]�j  K
j  KubK j  )��}�(h�jP  j  ]�j  K
j  K ubK!j  )��}�(h�jP  j  ]�j  K
j  K!ubK"j  )��}�(h�jP  j  ]�j  K
j  K"ubK#j  )��}�(h�jP  j  ]�j  K
j  K#ubK$j  )��}�(h�jP  j  ]�j  K
j  K$ubK%j  )��}�(h�jP  j  ]�j  K
j  K%ubK&j  )��}�(h�jP  j  ]�j  K
j  K&ubK'j  )��}�(h�jP  j  ]�j  K
j  K'ubK(j  )��}�(h�jP  j  ]�j  K
j  K(ubK)j  )��}�(h�jP  j  ]�j  K
j  K)ubK*j  )��}�(h�jP  j  ]�j  K
j  K*ubK+j  )��}�(h�jP  j  ]�j  K
j  K+ubK,j  )��}�(h�jP  j  ]�j  K
j  K,ubK-j  )��}�(h�jP  j  ]�j  K
j  K-ubK.j  )��}�(h�jP  j  ]�j  K
j  K.ubK/j  )��}�(h�jP  j  ]�j  K
j  K/ubK0j  )��}�(h�jP  j  ]�j  K
j  K0ubK1j  )��}�(h�jP  j  ]�j  K
j  K1ubK2j  )��}�(h�jP  j  ]�j  K
j  K2ubK3j  )��}�(h�jP  j  ]�j  K
j  K3ubK4j  )��}�(h�jP  j  ]�j  K
j  K4ubK5j  )��}�(h�jP  j  ]�j  K
j  K5ubK6j  )��}�(h�jP  j  ]�j  K
j  K6ubK7j  )��}�(h�jP  j  ]�j  K
j  K7ubK8j  )��}�(h�jP  j  ]�j  K
j  K8ubK9j  )��}�(h�jP  j  ]�j  K
j  K9ubK:j  )��}�(h�jP  j  ]�j  K
j  K:ubK;j  )��}�(h�jP  j  ]�j  K
j  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  �      ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�K
aj  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�Kaj  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�Kaj  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK}�(K j  )��}�(h�jP  j  ]�j  Kj  K ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK	j  )��}�(h�jP  j  ]�j  Kj  K	ubK
j  )��}�(h�jP  j  ]�j  Kj  K
ubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubKj  )��}�(h�jP  j  ]�j  Kj  KubK j  )��}�(h�jP  j  ]�j  Kj  K ubK!j  )��}�(h�jP  j  ]�j  Kj  K!ubK"j  )��}�(h�jP  j  ]�j  Kj  K"ubK#j  )��}�(h�jP  j  ]�j  Kj  K#ubK$j  )��}�(h�jP  j  ]�j  Kj  K$ubK%j  )��}�(h�jP  j  ]�j  Kj  K%ubK&j  )��}�(h�jP  j  ]�j  Kj  K&ubK'j  )��}�(h�jP  j  ]�j  Kj  K'ubK(j  )��}�(h�jP  j  ]�j  Kj  K(ubK)j  )��}�(h�jP  j  ]�j  Kj  K)ubK*j  )��}�(h�jP  j  ]�j  Kj  K*ubK+j  )��}�(h�jP  j  ]�j  Kj  K+ubK,j  )��}�(h�jP  j  ]�j  Kj  K,ubK-j  )��}�(h�jP  j  ]�j  Kj  K-ubK.j  )��}�(h�jP  j  ]�j  Kj  K.ubK/j  )��}�(h�jP  j  ]�j  Kj  K/ubK0j  )��}�(h�jP  j  ]�j  Kj  K0ubK1j  )��}�(h�jP  j  ]�j  Kj  K1ubK2j  )��}�(h�jP  j  ]�j  Kj  K2ubK3j  )��}�(h�jP  j  ]�j  Kj  K3ubK4j  )��}�(h�jP  j  ]�j  Kj  K4ubK5j  )��}�(h�jP  j  ]�j  Kj  K5ubK6j  )��}�(h�jP  j  ]�j  Kj  K6ubK7j  )��}�(h�jP  j  ]�j  Kj  K7ubK8j  )��}�(h�jP  j  ]�j  Kj  K8ubK9j  )��}�(h�jP  j  ]�j  Kj  K9ubK:j  )��}�(h�jP  j  ]�j  Kj  K:ubK;j  )��}�(h�jP  j  ]�j  Kj  K;ubuK }�(K j  )��}�(h�jP  j  ]�j  K j  K ubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubK	j  )��}�(h�jP  j  ]�j  K j  K	ubK
j  )��}�(h�jP  j  ]�j  K j  K
ubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubKj  )��}�(h�jP  j  ]�j  K j  KubK j  )��}�(h�jP  j  ]�j  K j  K ubK!j  )��}�(h�jP  j  ]�j  K j  K!ubK"j  )��}�(h�jP  j  ]�j  K j  K"ubK#j  )��}�(h�jP  j  ]�j  K j  K#ubK$j  )��}�(h�jP  j  ]�j  K j  K$ubK%j  )��}�(h�jP  j  ]�j  K j  K%ubK&j  )��}�(h�jP  j  ]�j  K j  K&ubK'j  )��}�(h�jP  j  ]�j  K j  K'ubK(j  )��}�(h�jP  j  ]�j  K j  K(ubK)j  )��}�(h�jP  j  ]�j  K j  K)ubK*j  )��}�(h�jP  j  ]�j  K j  K*ubK+j  )��}�(h�jP  j  ]�j  K j  K+ubK,j  )��}�(h�jP  j  ]�j  K j  K,ubK-j  )��}�(h�jP  j  ]�j  K j  K-ubK.j  )��}�(h�jP  j  ]�j  K j  K.ubK/j  )��}�(h�jP  j  ]�j  K j  K/ubK0j  )��}�(h�jP  j  ]�j  K j  K0ubK1j  )��}�(h�jP  j  ]�j  K j  K1ubK2j  )��}�(h�jP  j  ]�j  K j  K2ubK3j  )��}�(h�jP  j  ]�j  K j  K3ubK4j  )��}�(h�jP  j  ]�j  K j  K4ubK5j  )��}�(h�jP  j  ]�j  K j  K5ubK6j  )��}�(h�jP  j  ]�j  K j  K6ubK7j  )��}�(h�jP  j  ]�j  K j  K7ubK8j  )��}�(h�jP  j  ]�j  K j  K8ubK9j  )��}�(h�jP  j  ]�j  K j  K9ubK:j  )��}�(h�jP  j  ]�j  K j  K:ubK;j  )��}�(h�jP  j  ]�j  K j  K;ubuK!}�(K j  )��}�(h�jP  j  ]�j  K!j  K ubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubK	j  )��}�(h�jP  j  ]�j  K!j  K	ubK
j  )��}�(h�jP  j  ]�j  K!j  K
ubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubKj  )��}�(h�jP  j  ]�j  K!j  KubK j  )��}�(h�jP  j  ]�j  K!j  K ubK!j  )��}�(h�jP  j  ]�j  K!j  K!ubK"j  )��}�(h�jP  j  ]�j  K!j  K"ubK#j  )��}�(h�jP  j  ]�j  K!j  K#ubK$j  )��}�(h�jP  j  ]�j  K!j  K$ubK%j  )��}�(h�jP  j  ]�j  K!j  K%ubK&j  )��}�(h�jP  j  ]�j  K!j  K&ubK'j  )��}�(h�jP  j  ]�j  K!j  K'ubK(j  )��}�(h�jP  j  ]�j  K!j  K(ubK)j  )��}�(h�jP  j  ]�j  K!j  K)ubK*j  )��}�(h�jP  j  ]�j  K!j  K*ubK+j  )��}�(h�jP  j  ]�j  K!j  K+ubK,j  )��}�(h�jP  j  ]�j  K!j  K,ubK-j  )��}�(h�jP  j  ]�j  K!j  K-ubK.j  )��}�(h�jP  j  ]�j  K!j  K.ubK/j  )��}�(h�jP  j  ]�j  K!j  K/ubK0j  )��}�(h�jP  j  ]�j  K!j  K0ubK1j  )��}�(h�jP  j  ]�j  K!j  K1ubK2j  )��}�(h�jP  j  ]�j  K!j  K2ubK3j  )��}�(h�jP  j  ]�j  K!j  K3ubK4j  )��}�(h�jP  j  ]�j  K!j  K4ubK5j  )��}�(h�jP  j  ]�j  K!j  K5ubK6j  )��}�(h�jP  j  ]�j  K!j  K6ubK7j  )��}�(h�jP  j  ]�j  K!j  K7ubK8j  )��}�(h�jP  j  ]�j  K!j  K8ubK9j  )��}�(h�jP  j  ]�j  K!j  K9ubK:j  )��}�(h�jP  j  ]�j  K!j  K:ubK;j  )��}�(h�jP  j  ]�j  K!j  K;ubuK"}�(K j  )��}�(h�jP  j  ]�j  K"j  K ubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubK	j  )��}�(h�jP  j  ]�j  K"j  K	ubK
j  )��}�(h�jP  j  ]�j  K"j  K
ubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubKj  )��}�(h�jP  j  ]�j  K"j  KubK j  )��}�(h�jP  j  ]�j  K"j  K ubK!j  )��}�(h�jP  j  ]�j  K"j  K!ubK"j  )��}�(h�jP  j  ]�j  K"j  K"ubK#j  )��}�(h�jP  j  ]�j  K"j  K#ubK$j  )��}�(h�jP  j  ]�j  K"j  K$ubK%j  )��}�(h�jP  j  ]�j  K"j  K%ubK&j  )��}�(h�jP  j  ]�j  K"j  K&ubK'j  )��}�(h�jP  j  ]�j  K"j  K'ubK(j  )��}�(h�jP  j  ]�j  K"j  K(ubK)j  )��}�(h�jP  j  ]�j  K"j  K)ubK*j  )��}�(h�jP  j  ]�j  K"j  K*ubK+j  )��}�(h�jP  j  ]�j  K"j  K+ubK,j  )��}�(h�jP  j  ]�j  K"j  K,ubK-j  )��}�(h�jP  j  ]�j  K"j  K-ubK.j  )��}�(h�jP  j  ]�j  K"j  K.ubK/j  )��}�(h�jP  j  ]�j  K"j  K/ubK0j  )��}�(h�jP  j  ]�j  K"j  K0ubK1j  )��}�(h�jP  j  ]�j  K"j  K1ubK2j  )��}�(h�jP  j  ]�j  K"j  K2ubK3j  )��}�(h�jP  j  ]�j  K"j  K3ubK4j  )��}�(h�jP  j  ]�j  K"j  K4ubK5j  )��}�(h�jP  j  ]�j  K"j  K5ubK6j  )��}�(h�jP  j  ]�j  K"j  K6ubK7j  )��}�(h�jP  j  ]�j  K"j  K7ubK8j  )��}�(h�jP  j  ]�j  K"j  K8ubK9j  )��}�(h�jP  j  ]�j  K"j  K9ubK:j  )��}�(h�jP  j  ]�j  K"j  K:ubK;j  )��}�(h�jP  j  ]�j  K"j  K;ubuK#}�(K j  )��}�(h�jP  j  ]�j  K#j  K ubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubK	j  )��}�(h�jP  j  ]�j  K#j  K	ubK
j  )��}�(h�jP  j  ]�j  K#j  K
ubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubKj  )��}�(h�jP  j  ]�j  K#j  KubK j  )��}�(h�jP  j  ]�j  K#j  K ubK!j  )��}�(h�jP  j  ]�j  K#j  K!ubK"j  )��}�(h�jP  j  ]�j  K#j  K"ubK#j  )��}�(h�jP  j  ]�j  K#j  K#ubK$j  )��}�(h�jP  j  ]�j  K#j  K$ubK%j  )��}�(h�jP  j  ]�j  K#j  K%ubK&j  )��}�(h�jP  j  ]�j  K#j  K&ubK'j  )��}�(h�jP  j  ]�j  K#j  K'ubK(j  )��}�(h�jP  j  ]�j  K#j  K(ubK)j  )��}�(h�jP  j  ]�j  K#j  K)ubK*j  )��}�(h�jP  j  ]�j  K#j  K*ubK+j  )��}�(h�jP  j  ]�j  K#j  K+ubK,j  )��}�(h�jP  j  ]�j  K#j  K,ubK-j  )��}�(h�jP  j  ]�j  K#j  K-ubK.j  )��}�(h�jP  j  ]�j  K#j  K.ubK/j  )��}�(h�jP  j  ]�j  K#j  K/ubK0j  )��}�(h�jP  j  ]�j  K#j  K0ubK1j  )��}�(h�jP  j  ]�j  K#j  K1ubK2j  )��}�(h�jP  j  ]�j  K#j  K2ubK3j  )��}�(h�jP  j  ]�j  K#j  K3ubK4j  )��}�(h�jP  j  ]�j  K#j  K4ubK5j  )��}�(h�jP  j  ]�j  K#j  K5ubK6j  )��}�(h�jP  j  ]�j  K#j  K6ubK7j  )��}�(h�jP  j  ]�j  K#j  K7ubK8j  )��}�(h�jP  j  ]�j  K#j  K8ubK9j  )��}�(h�jP  j  ]�j  K#j  K9ubK:j  )��}�(h�jP  j  ]�j  K#j  K:ubK;j  )��}�(h�jP  j  ]�j  K#j  K;ubuK$}�(K j  )��}�(h�jP  j  ]�j  K$j  K ubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubK	j  )��}�(h�jP  j  ]�j  K$j  K	ubK
j  )��}�(h�jP  j  ]�j  K$j  K
ubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubKj  )��}�(h�jP  j  ]�j  K$j  KubK j  )��}�(h�jP  j  ]�j  K$j  K ubK!j  )��}�(h�jP  j  ]�j  K$j  K!ubK"j  )��}�(h�jP  j  ]�j  K$j  K"ubK#j  )��}�(h�jP  j  ]�j  K$j  K#ubK$j  )��}�(h�jP  j  ]�j  K$j  K$ubK%j  )��}�(h�jP  j  ]�j  K$j  K%ubK&j  )��}�(h�jP  j  ]�j  K$j  K&ubK'j  )��}�(h�jP  j  ]�j  K$j  K'ubK(j  )��}�(h�jP  j  ]�j  K$j  K(ubK)j  )��}�(h�jP  j  ]�j  K$j  K)ubK*j  )��}�(h�jP  j  ]�j  K$j  K*ubK+j  )��}�(h�jP  j  ]�j  K$j  K+ubK,j  )��}�(h�jP  j  ]�j  K$j  K,ubK-j  )��}�(h�jP  j  ]�j  K$j  K-ubK.j  )��}�(h�jP  j  ]�j  K$j  K.ubK/j  )��}�(h�jP  j  ]�j  K$j  K/ubK0j  )��}�(h�jP  j  ]�j  K$j  K0ubK1j  )��}�(h�jP  j  ]�j  K$j  K1ubK2j  )��}�(h�jP  j  ]�j  K$j  K2ubK3j  )��}�(h�jP  j  ]�j  K$j  K3ubK4j  )��}�(h�jP  j  ]�j  K$j  K4ubK5j  )��}�(h�jP  j  ]�j  K$j  K5ubK6j  )��}�(h�jP  j  ]�j  K$j  K6ubK7j  )��}�(h�jP  j  ]�j  K$j  K7ubK8j  )��}�(h�jP  j  ]�j  K$j  K8ubK9j  )��}�(h�jP  j  ]�j  K$j  K9ubK:j  )��}�(h�jP  j  ]�j  K$j  K:ubK;j  )��}�(h�jP  j  ]�j  K$j  K;ubuK%}�(K j  )��}�(h�jP  j  ]�j  K%j  K ubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubK	j  )��}�(h�jP  j  ]�j  K%j  K	ubK
j  )��}�(h�jP  j  ]�j  K%j  K
ubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubKj  )��}�(h�jP  j  ]�j  K%j  KubK j  )��}�(h�jP  j  ]�j  K%j  K ubK!j  )��}�(h�jP  j  ]�j  K%j  K!ubK"j  )��}�(h�jP  j  ]�j  K%j  K"ubK#j  )��}�(h�jP  j  ]�j  K%j  K#ubK$j  )��}�(h�jP  j  ]�j  K%j  K$ubK%j  )��}�(h�jP  j  ]�j  K%j  K%ub�       K&j  )��}�(h�jP  j  ]�j  K%j  K&ubK'j  )��}�(h�jP  j  ]�j  K%j  K'ubK(j  )��}�(h�jP  j  ]�j  K%j  K(ubK)j  )��}�(h�jP  j  ]�j  K%j  K)ubK*j  )��}�(h�jP  j  ]�j  K%j  K*ubK+j  )��}�(h�jP  j  ]�j  K%j  K+ubK,j  )��}�(h�jP  j  ]�j  K%j  K,ubK-j  )��}�(h�jP  j  ]�j  K%j  K-ubK.j  )��}�(h�jP  j  ]�j  K%j  K.ubK/j  )��}�(h�jP  j  ]�j  K%j  K/ubK0j  )��}�(h�jP  j  ]�j  K%j  K0ubK1j  )��}�(h�jP  j  ]�j  K%j  K1ubK2j  )��}�(h�jP  j  ]�j  K%j  K2ubK3j  )��}�(h�jP  j  ]�j  K%j  K3ubK4j  )��}�(h�jP  j  ]�j  K%j  K4ubK5j  )��}�(h�jP  j  ]�j  K%j  K5ubK6j  )��}�(h�jP  j  ]�j  K%j  K6ubK7j  )��}�(h�jP  j  ]�j  K%j  K7ubK8j  )��}�(h�jP  j  ]�j  K%j  K8ubK9j  )��}�(h�jP  j  ]�j  K%j  K9ubK:j  )��}�(h�jP  j  ]�j  K%j  K:ubK;j  )��}�(h�jP  j  ]�j  K%j  K;ubuK&}�(K j  )��}�(h�jP  j  ]�j  K&j  K ubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubK	j  )��}�(h�jP  j  ]�j  K&j  K	ubK
j  )��}�(h�jP  j  ]�j  K&j  K
ubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubKj  )��}�(h�jP  j  ]�j  K&j  KubK j  )��}�(h�jP  j  ]�j  K&j  K ubK!j  )��}�(h�jP  j  ]�j  K&j  K!ubK"j  )��}�(h�jP  j  ]�j  K&j  K"ubK#j  )��}�(h�jP  j  ]�j  K&j  K#ubK$j  )��}�(h�jP  j  ]�j  K&j  K$ubK%j  )��}�(h�jP  j  ]�j  K&j  K%ubK&j  )��}�(h�jP  j  ]�j  K&j  K&ubK'j  )��}�(h�jP  j  ]�j  K&j  K'ubK(j  )��}�(h�jP  j  ]�j  K&j  K(ubK)j  )��}�(h�jP  j  ]�j  K&j  K)ubK*j  )��}�(h�jP  j  ]�j  K&j  K*ubK+j  )��}�(h�jP  j  ]�j  K&j  K+ubK,j  )��}�(h�jP  j  ]�j  K&j  K,ubK-j  )��}�(h�jP  j  ]�j  K&j  K-ubK.j  )��}�(h�jP  j  ]�j  K&j  K.ubK/j  )��}�(h�jP  j  ]�j  K&j  K/ubK0j  )��}�(h�jP  j  ]�j  K&j  K0ubK1j  )��}�(h�jP  j  ]�j  K&j  K1ubK2j  )��}�(h�jP  j  ]�j  K&j  K2ubK3j  )��}�(h�jP  j  ]�j  K&j  K3ubK4j  )��}�(h�jP  j  ]�j  K&j  K4ubK5j  )��}�(h�jP  j  ]�j  K&j  K5ubK6j  )��}�(h�jP  j  ]�j  K&j  K6ubK7j  )��}�(h�jP  j  ]�j  K&j  K7ubK8j  )��}�(h�jP  j  ]�j  K&j  K8ubK9j  )��}�(h�jP  j  ]�j  K&j  K9ubK:j  )��}�(h�jP  j  ]�j  K&j  K:ubK;j  )��}�(h�jP  j  ]�j  K&j  K;ubuK'}�(K j  )��}�(h�jP  j  ]�j  K'j  K ubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubK	j  )��}�(h�jP  j  ]�j  K'j  K	ubK
j  )��}�(h�jP  j  ]�j  K'j  K
ubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubKj  )��}�(h�jP  j  ]�j  K'j  KubK j  )��}�(h�jP  j  ]�j  K'j  K ubK!j  )��}�(h�jP  j  ]�j  K'j  K!ubK"j  )��}�(h�jP  j  ]�j  K'j  K"ubK#j  )��}�(h�jP  j  ]�j  K'j  K#ubK$j  )��}�(h�jP  j  ]�j  K'j  K$ubK%j  )��}�(h�jP  j  ]�j  K'j  K%ubK&j  )��}�(h�jP  j  ]�j  K'j  K&ubK'j  )��}�(h�jP  j  ]�j  K'j  K'ubK(j  )��}�(h�jP  j  ]�j  K'j  K(ubK)j  )��}�(h�jP  j  ]�j  K'j  K)ubK*j  )��}�(h�jP  j  ]�j  K'j  K*ubK+j  )��}�(h�jP  j  ]�j  K'j  K+ubK,j  )��}�(h�jP  j  ]�j  K'j  K,ubK-j  )��}�(h�jP  j  ]�j  K'j  K-ubK.j  )��}�(h�jP  j  ]�j  K'j  K.ubK/j  )��}�(h�jP  j  ]�j  K'j  K/ubK0j  )��}�(h�jP  j  ]�j  K'j  K0ubK1j  )��}�(h�jP  j  ]�j  K'j  K1ubK2j  )��}�(h�jP  j  ]�j  K'j  K2ubK3j  )��}�(h�jP  j  ]�j  K'j  K3ubK4j  )��}�(h�jP  j  ]�j  K'j  K4ubK5j  )��}�(h�jP  j  ]�j  K'j  K5ubK6j  )��}�(h�jP  j  ]�j  K'j  K6ubK7j  )��}�(h�jP  j  ]�j  K'j  K7ubK8j  )��}�(h�jP  j  ]�j  K'j  K8ubK9j  )��}�(h�jP  j  ]�j  K'j  K9ubK:j  )��}�(h�jP  j  ]�j  K'j  K:ubK;j  )��}�(h�jP  j  ]�j  K'j  K;ubuK(}�(K j  )��}�(h�jP  j  ]�j  K(j  K ubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubK	j  )��}�(h�jP  j  ]�j  K(j  K	ubK
j  )��}�(h�jP  j  ]�j  K(j  K
ubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubKj  )��}�(h�jP  j  ]�j  K(j  KubK j  )��}�(h�jP  j  ]�j  K(j  K ubK!j  )��}�(h�jP  j  ]�j  K(j  K!ubK"j  )��}�(h�jP  j  ]�j  K(j  K"ubK#j  )��}�(h�jP  j  ]�j  K(j  K#ubK$j  )��}�(h�jP  j  ]�j  K(j  K$ubK%j  )��}�(h�jP  j  ]�Kaj  K(j  K%ubK&j  )��}�(h�jP  j  ]�j  K(j  K&ubK'j  )��}�(h�jP  j  ]�j  K(j  K'ubK(j  )��}�(h�jP  j  ]�j  K(j  K(ubK)j  )��}�(h�jP  j  ]�(KKej  K(j  K)ubK*j  )��}�(h�jP  j  ]�j  K(j  K*ubK+j  )��}�(h�jP  j  ]�j  K(j  K+ubK,j  )��}�(h�jP  j  ]�j  K(j  K,ubK-j  )��}�(h�jP  j  ]�j  K(j  K-ubK.j  )��}�(h�jP  j  ]�j  K(j  K.ubK/j  )��}�(h�jP  j  ]�j  K(j  K/ubK0j  )��}�(h�jP  j  ]�j  K(j  K0ubK1j  )��}�(h�jP  j  ]�j  K(j  K1ubK2j  )��}�(h�jP  j  ]�j  K(j  K2ubK3j  )��}�(h�jP  j  ]�j  K(j  K3ubK4j  )��}�(h�jP  j  ]�j  K(j  K4ubK5j  )��}�(h�jP  j  ]�j  K(j  K5ubK6j  )��}�(h�jP  j  ]�j  K(j  K6ubK7j  )��}�(h�jP  j  ]�j  K(j  K7ubK8j  )��}�(h�jP  j  ]�j  K(j  K8ubK9j  )��}�(h�jP  j  ]�j  K(j  K9ubK:j  )��}�(h�jP  j  ]�j  K(j  K:ubK;j  )��}�(h�jP  j  ]�j  K(j  K;ubuK)}�(K j  )��}�(h�jP  j  ]�j  K)j  K ubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubK	j  )��}�(h�jP  j  ]�j  K)j  K	ubK
j  )��}�(h�jP  j  ]�j  K)j  K
ubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubKj  )��}�(h�jP  j  ]�j  K)j  KubK j  )��}�(h�jP  j  ]�j  K)j  K ubK!j  )��}�(h�jP  j  ]�j  K)j  K!ubK"j  )��}�(h�jP  j  ]�j  K)j  K"ubK#j  )��}�(h�jP  j  ]�j  K)j  K#ubK$j  )��}�(h�jP  j  ]�j  K)j  K$ubK%j  )��}�(h�jP  j  ]�j  K)j  K%ubK&j  )��}�(h�jP  j  ]�j  K)j  K&ubK'j  )��}�(h�jP  j  ]�Kaj  K)j  K'ubK(j  )��}�(h�jP  j  ]�j  K)j  K(ubK)j  )��}�(h�jP  j  ]�j  K)j  K)ubK*j  )��}�(h�jP  j  ]�j  K)j  K*ubK+j  )��}�(h�jP  j  ]�j  K)j  K+ubK,j  )��}�(h�jP  j  ]�j  K)j  K,ubK-j  )��}�(h�jP  j  ]�j  K)j  K-ubK.j  )��}�(h�jP  j  ]�j  K)j  K.ubK/j  )��}�(h�jP  j  ]�j  K)j  K/ubK0j  )��}�(h�jP  j  ]�j  K)j  K0ubK1j  )��}�(h�jP  j  ]�j  K)j  K1ubK2j  )��}�(h�jP  j  ]�j  K)j  K2ubK3j  )��}�(h�jP  j  ]�j  K)j  K3ubK4j  )��}�(h�jP  j  ]�j  K)j  K4ubK5j  )��}�(h�jP  j  ]�j  K)j  K5ubK6j  )��}�(h�jP  j  ]�j  K)j  K6ubK7j  )��}�(h�jP  j  ]�j  K)j  K7ubK8j  )��}�(h�jP  j  ]�j  K)j  K8ubK9j  )��}�(h�jP  j  ]�j  K)j  K9ubK:j  )��}�(h�jP  j  ]�j  K)j  K:ubK;j  )��}�(h�jP  j  ]�j  K)j  K;ubuK*}�(K j  )��}�(h�jP  j  ]�j  K*j  K ubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubK	j  )��}�(h�jP  j  ]�j  K*j  K	ubK
j  )��}�(h�jP  j  ]�j  K*j  K
ubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubKj  )��}�(h�jP  j  ]�j  K*j  KubK j  )��}�(h�jP  j  ]�j  K*j  K ubK!j  )��}�(h�jP  j  ]�j  K*j  K!ubK"j  )��}�(h�jP  j  ]�j  K*j  K"ubK#j  )��}�(h�jP  j  ]�j  K*j  K#ubK$j  )��}�(h�jP  j  ]�j  K*j  K$ubK%j  )��}�(h�jP  j  ]�j  K*j  K%ubK&j  )��}�(h�jP  j  ]�j  K*j  K&ubK'j  )��}�(h�jP  j  ]�j  K*j  K'ubK(j  )��}�(h�jP  j  ]�j  K*j  K(ubK)j  )��}�(h�jP  j  ]�j  K*j  K)ubK*j  )��}�(h�jP  j  ]�j  K*j  K*ubK+j  )��}�(h�jP  j  ]�j  K*j  K+ubK,j  )��}�(h�jP  j  ]�j  K*j  K,ubK-j  )��}�(h�jP  j  ]�j  K*j  K-ubK.j  )��}�(h�jP  j  ]�j  K*j  K.ubK/j  )��}�(h�jP  j  ]�j  K*j  K/ubK0j  )��}�(h�jP  j  ]�j  K*j  K0ubK1j  )��}�(h�jP  j  ]�j  K*j  K1ubK2j  )��}�(h�jP  j  ]�j  K*j  K2ubK3j  )��}�(h�jP  j  ]�j  K*j  K3ubK4j  )��}�(h�jP  j  ]�j  K*j  K4ubK5j  )��}�(h�jP  j  ]�j  K*j  K5ubK6j  )��}�(h�jP  j  ]�j  K*j  K6ubK7j  )��}�(h�jP  j  ]�j  K*j  K7ubK8j  )��}�(h�jP  j  ]�j  K*j  K8ubK9j  )��}�(h�jP  j  ]�j  K*j  K9ubK:j  )��}�(h�jP  j  ]�j  K*j  K:ubK;j  )��}�(h�jP  j  ]�j  K*j  K;ubuK+}�(K j  )��}�(h�jP  j  ]�j  K+j  K ubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubK	j  )��}�(h�jP  j  ]�j  K+j  K	ubK
j  )��}�(h�jP  j  ]�j  K+j  K
ubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubKj  )��}�(h�jP  j  ]�j  K+j  KubK j  )��}�(h�jP  j  ]�j  K+j  K ubK!j  )��}�(h�jP  j  ]�j  K+j  K!ubK"j  )��}�(h�jP  j  ]�j  K+j  K"ubK#j  )��}�(h�jP  j  ]�j  K+j  K#ubK$j  )��}�(h�jP  j  ]�j  K+j  K$ubK%j  )��}�(h�jP  j  ]�j  K+j  K%ubK&j  )��}�(h�jP  j  ]�j  K+j  K&ubK'j  )��}�(h�jP  j  ]�j  K+j  K'ubK(j  )��}�(h�jP  j  ]�j  K+j  K(ubK)j  )��}�(h�jP  j  ]�j  K+j  K)ubK*j  )��}�(h�jP  j  ]�j  K+j  K*ubK+j  )��}�(h�jP  j  ]�j  K+j  K+ubK,j  )��}�(h�jP  j  ]�j  K+j  K,ubK-j  )��}�(h�jP  j  ]�j  K+j  K-ubK.j  )��}�(h�jP  j  ]�j  K+j  K.ubK/j  )��}�(h�jP  j  ]�j  K+j  K/ubK0j  )��}�(h�jP  j  ]�j  K+j  K0ubK1j  )��}�(h�jP  j  ]�j  K+j  K1ubK2j  )��}�(h�jP  j  ]�j  K+j  K2ubK3j  )��}�(h�jP  j  ]�j  K+j  K3ubK4j  )��}�(h�jP  j  ]�j  K+j  K4ubK5j  )��}�(h�jP  j  ]�j  K+j  K5ubK6j  )��}�(h�jP  j  ]�j  K+j  K6ubK7j  )��}�(h�jP  j  ]�j  K+j  K7ubK8j  )��}�(h�jP  j  ]�j  K+j  K8ubK9j  )��}�(h�jP  j  ]�j  K+j  K9ubK:j  )��}�(h�jP  j  ]�j  K+j  K:ubK;j  )��}�(h�jP  j  ]�j  K+j  K;ubuK,}�(K j  )��}�(h�jP  j  ]�j  K,j  K ubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubK	j  )��}�(h�jP  j  ]�j  K,j  K	ubK
j  )��}�(h�jP  j  ]�j  K,j  K
ubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubKj  )��}�(h�jP  j  ]�j  K,j  KubK j  )��}�(h�jP  j  ]�j  K,j  K ubK!j  )��}�(h�jP  j  ]�j  K,j  K!ubK"j  )��}�(h�jP  j  ]�j  K,j  K"ubK#j  )��}�(h�jP  j  ]�j  K,j  K#ubK$j  )��}�(h�jP  j  ]�j  K,j  K$ubK%j  )��}�(h�jP  j  ]�j  K,j  K%ubK&j  )��}�(h�jP  j  ]�j  K,j  K&ubK'j  )��}�(h�jP  j  ]�j  K,j  K'ubK(j  )��}�(h�jP  j  ]�j  K,j  K(ubK)j  )��}�(h�jP  j  ]�j  K,j  K)ubK*j  )��}�(h�jP  j  ]�j  K,j  K*ubK+j  )��}�(h�jP  j  ]�j  K,j  K+ubK,j  )��}�(h�jP  j  ]�j  K,j  K,ubK-j  )��}�(h�jP  j  ]�j  K,j  K-ubK.j  )��}�(h�jP  j  ]�j  K,j  K.ubK/j  )��}�(h�jP  j  ]�j  K,j  K/ubK0j  )��}�(h�jP  j  ]�j  K,j  K0ubK1j  )��}�(h�jP  j  ]�j  K,j  K1ubK2j  )��}�(h�jP  j  ]�j  K,j  K2ubK3j  )��}�(h�jP  j  ]�j  K,j  K3ubK4j  )��}�(h�jP  j  ]�j  K,j  K4ubK5j  )��}�(h�jP  j  ]�j  K,j  K5ubK6j  )��}�(h�jP  j  ]�j  K,j  K6ubK7j  )��}�(h�jP  j  ]�j  K,j  K7ubK8j  )��}�(h�jP  j  ]�j  K,j  K8ubK9j  )��}�(h�jP  j  ]�j  K,j  K9ubK:j  )��}�(h�jP  j  ]�j  K,j  K:ubK;j  )��}�(h�jP  j  ]�j  K,j  K;ubuK-}�(K j  )��}�(h�jP  j  ]�j  K-j  K ubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubK	j  )��}�(h�jP  j  ]�j  K-j  K	ubK
j  )��}�(h�jP  j  ]�j  K-j  K
ubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubKj  )��}�(h�jP  j  ]�j  K-j  KubK j  )��}�(h�jP  j  ]�j  K-j  K ubK!j  )��}�(h�jP  j  ]�j  K-j  K!ubK"j  )��}�(h�jP  j  ]�j  K-j  K"ubK#j  )��}�(h�jP  j  ]�j  K-j  K#ubK$j  )��}�(h�jP  j  ]�j  K-j  K$ubK%j  )��}�(h�jP  j  ]�Kaj  K-j  K%ubK&j  )��}�(h�jP  j  ]�j  K-j  K&ubK'j  )��}�(h�jP  j  ]�j  K-j  K'ubK(j  )��}�(h�jP  j  ]�j  K-j  K(ubK)j  )��}�(h�jP  j  ]�j  K-j  K)ubK*j  )��}�(h�jP  j  ]�j  K-j  K*ubK+j  )��}�(h�jP  j  ]�j  K-j  K+ubK,j  )��}�(h�jP  j  ]�j  K-j  K,ubK-j  )��}�(h�jP  j  ]�j  K-j  K-ubK.j  )��}�(h�jP  j  ]�j  K-j  K.ubK/j  )��}�(h�jP  j  ]�j  K-j  K/ubK0j  )��}�(h�jP  j  ]�j  K-j  K0ubK1j  )��}�(h�jP  j  ]�j  K-j  K1ubK2j  )��}�(h�jP  j  ]�j  K-j  K2ubK3j  )��}�(h�jP  j  ]�j  K-j  K3ubK4j  )��}�(h�jP  j  ]�j  K-j  K4ubK5j  )��}�(h�jP  j  ]�j  K-j  K5ubK6j  )��}�(h�jP  j  ]�j  K-j  K6ubK7j  )��}�(h�jP  j  ]�j  K-j  K7ubK8j  )��}�(h�jP  j  ]�j  K-j  K8ubK9j  )��}�(h�jP  j  ]�j  K-j  K9ubK:j  )��}�(h�jP  j  ]�j  K-j  K:ubK;j  )��}�(h�jP  j  ]�j  K-j  K;ubuK.}�(K j  )��}�(h�jP  j  ]�j  K.j  K ubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubK	j  )��}�(h�jP  j  ]�j  K.j  K	ubK
j  )��}�(h�jP  j  ]�j  K.j  K
ubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubKj  )��}�(h�jP  j  ]�j  K.j  KubK j  )��}�(h�jP  j  ]�j  K.j  K ubK!j  )��}�(h�jP  j  ]�j  K.j  K!ubK"j  )��}�(h�jP  j  ]�j  K.j  K"ubK#j  )��}�(h�jP  j  ]�j  K.j  K#ubK$j  )��}�(h�jP  j  ]�j  K.j  K$ubK%j  )��}�(h�jP  j  ]�j  K.j  K%ubK&j  )��}�(h�jP  j  ]�j  K.j  K&ubK'j  )��}�(h�jP  j  ]�j  K.j  K'ubK(j  )��}�(h�jP  j  ]�j  K.j  K(ubK)j  )��}�(h�jP  j  ]�j  K.j  K)ubK*j  )��}�(h�jP  j  ]�j  K.j  K*ubK+j  )��}�(h�jP  j  ]�j  K.j  K+ubK,j  )��}�(h�jP  j  ]�j  K.j  K,ubK-j  )��}�(h�jP  j  ]�j  K.j  K-ubK.j  )��}�(h�jP  j  ]�j  K.j  K.ubK/j  )��}�(h�jP  j  ]�j  K.j  K/ubK0j  )��}�(h�jP  j  ]�j  K.j  K0ubK1j  )��}�(h�jP  j  ]�j  K.j  K1ubK2j  )��}�(h�jP  j  ]�j  K.j  K2ubK3j  )��}�(h�jP  j  ]�j  K.j  K3ubK4j  )��}�(h�jP  j  ]�j  K.j  K4ubK5j  )��}�(h�jP  j  ]�j  K.j  K5ubK6j  )��}�(h�jP  j  ]�j  K.j  K6ubK7j  )��}�(h�jP  j  ]�j  K.j  K7ubK8j  )��}�(h�jP  j  ]�j  K.j  K8ubK9j  )��}�(h�jP  j  ]�j  K.j  K9ubK:j  )��}�(h�jP  j  ]�j  K.j  K:ubK;j  )��}�(h�jP  j  ]�j  K.j  K;ubuK/}�(K j  )��}�(h�jP  j  ]�j  K/j  K ubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubK	j  )��}�(h�jP  j  ]�j  K/j  K	ubK
j  )��}�(h�jP  j  ]�j  K/j  K
ubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubKj  )��}�(h�jP  j  ]�j  K/j  KubK j  )��}�(h�jP  j  ]�j  K/j  K ubK!j  )��}�(h�jP  j  ]�j  K/j  K!ubK"j  )��}�(h�jP  j  ]�j  K/j  K"ubK#j  )��}�(h�jP  j  ]�j  K/j  K#ubK$j  )��}�(h�jP  j  ]�j  K/j  K$ubK%j  )��}�(h�jP  j  ]�j  K/j  K%ubK&j  )��}�(h�jP  j  ]�j  K/j  K&ubK'j  )��}�(h�jP  j  ]�j  K/j  K'ubK(j  )��}�(h�jP  j  ]�j  K/j  K(ubK)j  )��}�(h�jP  j  ]�j  K/j  K)ubK*j  )��}�(h�jP  j  ]�j  K/j  K*ubK+j  )��}�(h�jP  j  ]�j  K/j  K+ubK,j  )��}�(h�jP  j  ]�j  K/j  K,ubK-j  )��}�(h�jP  j  ]�j  K/j  K-ubK.j  )��}�(h�jP  j  ]�j  K/j  K.ubK/j  )��}�(h�jP  j  ]�j  K/j  K/ubK0j  )��}�(h�jP  j  ]�j  K/j  K0ubK1j  )��}�(h�jP  j  ]�j  K/j  K1ubK2j  )��}�(h�jP  j  ]�j  K/j  K2ubK3j  )��}�(h�jP  j  ]�j  K/j  K3ubK4j  )��}�(h�jP  j  ]�j  K/j  K4ubK5j  )��}�(h�jP  j  ]�j  K/j  K5ubK6j  )��}�(h�jP  j  ]�j  K/j  K6ubK7j  )��}�(h�jP  j  ]�j  K/j  K7ubK8j  )��}�(h�jP  j  ]�j  K/j  K8ubK9j  )��}�(h�jP  j  ]�j  K/j  K9ubK:j  )��}�(h�jP  j  ]�j  K/j  K:ubK;j  )��}�(h�jP  j  ]�j  K/j  K;ubuK0}�(K j  )��}�(h�jP  j  ]�j  K0j  K ubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubK	j  )��}�(h�jP  j  ]�j  K0j  K	ubK
j  )��}�(h�jP  j  ]�j  K0j  K
ubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubKj  )��}�(h�jP  j  ]�j  K0j  KubK j  )��}�(h�jP  j  ]�j  K0j  K ubK!j  )��}�(h�jP  j  ]�j  K0j  K!ubK"j  )��}�(h�jP  j  ]�j  K0j  K"ubK#j  )��}�(h�jP  j  ]�j  K0j  K#ubK$j  )��}�(h�jP  j  ]�j  K0j  K$ubK%j  )��}�(h�jP  j  ]�j  K0j  K%ubK&j  )��}�(h�jP  j  ]�j  K0j  K&ubK'j  )��}�(h�jP  j  ]�j  K0j  K'ubK(j  )��}�(h�jP  j  ]�j  K0j  K(ubK)j  )��}�(h�jP  j  ]�j  K0j  K)ubK*j  )��}�(h�jP  j  ]�j  K0j  K*ubK+j  )��}�(h�jP  j  ]�j  K0j  K+ubK,j  )��}�(h�jP  j  ]�j  K0j  K,ubK-j  )��}�(h�jP  j  ]�j  K0j  K-ubK.j  )��}�(h�jP  j  ]�j  K0j  K.ubK/j  )��}�(h�jP  j  ]�j  K0j  K/ubK0j  )��}�(h�jP  j  ]�j  K0j  K0ubK1j  )��}�(h�jP  j  ]�j  K0j  K1ubK2j  )��}�(h�jP  j  ]�j  K0j  K2ubK3j  )��}�(h�jP  j  ]�j  K0j  K3ubK4j  )��}�(h�jP  j  ]�j  K0j  K4ubK5j  )��}�(h�jP  j  ]�j  K0j  K5ubK6j  )��}�(h�jP  j  ]�j  K0j  K6ubK7j  )��}�(h�jP  j  ]�j  K0j  K7ubK8j  )��}�(h�jP  j  ]�j  K0j  K8ubK9j  )��}�(h�jP  j  ]�j  K0j  K9ubK:j  )��}�(h�jP  j  ]�j  K0j  K:ubK;j  )��}�(h�jP  j  ]�j  K0j  K;ubuK1}�(K j  )��}�(h�jP  j  ]�j  K1j  K ubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubK	j  )��}�(h�jP  j  ]�j  K1j  K	ubK
j  )��}�(h�jP  j  ]�j  K1j  K
ubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubKj  )��}�(h�jP  j  ]�j  K1j  KubK j  )��}�(h�jP  j  ]�j  K1j  K ubK!j  )��}�(h�jP  j  ]�j  K1j  K!ubK"j  )��}�(h�jP  j  ]�j  K1j  K"ubK#j  )��}�(h�jP  j  ]�j  K1j  K#ubK$j  )��}�(h�jP  j  ]�j  K1j  K$ubK%j  )��}�(h�jP  j  ]�j  K1j  K%ubK&j  )��}�(h�jP  j  ]�j  K1j  K&ubK'j  )��}�(h�jP  j  ]�j  K1j  K'ubK(j  )��}�(h�jP  j  ]�j  K1j  K(ubK)j  )��}�(h�jP  j  ]�j  K1j  K)ubK*j  )��}�(h�jP  j  ]�j  K1j  K*ubK+j  )��}�(h�jP  j  ]�j  K1j  K+ubK,j  )��}�(h�jP  j  ]�j  K1j  K,ubK-j  )��}�(h�jP  j  ]�j  K1j  K-ubK.j  )��}�(h�jP  j  ]�j  K1j  K.ubK/j  )��}�(h�jP  j  ]�j  K1j  K/ubK0j  )��}�(h�jP  j  ]�j  K1j  K0ubK1j  )��}�(h�jP  j  ]�j  K1j  K1ubK2j  )��}�(h�jP  j  ]�j  K1j  K2ubK3j  )��}�(h�jP  j  ]�j  K1j  K3ubK4j  )��}�(h�jP  j  ]�j  K1j  K4ubK5j  )��}�(h�jP  j  ]�j  K1j  K5ubK6j  )��}�(h�jP  j  ]�j  K1j  K6ubK7j  )��}�(h�jP  j  ]�j  K1j  K7ubK8j  )��}�(h�jP  j  ]�j  K1j  K8ubK9j  )��}�(h�jP  j  ]�j  K1j  K9ubK:j  )��}�(h�jP  j  ]�j  K1j  K:ubK;j  )��}�(h�jP  j  ]�j  K1j  K;ubuK2}�(K j  )��}�(h�jP  j  ]�j  K2j  K ubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubK	j  )��}�(h�jP  j  ]�j  K2j  K	ubK
j  )��}�(h�jP  j  ]�j  K2j  K
ubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubKj  )��}�(h�jP  j  ]�j  K2j  KubK j  )��}�(h�jP  j  ]�j  K2j  K ubK!j  )��}�(h�jP  j  ]�j  K2j  K!ubK"j  )��}�(h�jP  j  ]�j  K2j  K"ubK#j  )��}�(h�jP  j  ]�j  K2j  K#ubK$j  )��}�(h�jP  j  ]�j  K2j  K$ubK%j  )��}�(h�jP  j  ]�j  K2j  K%ubK&j  )��}�(h�jP  j  ]�j  K2j  K&ubK'j  )��}�(h�jP  j  ]�j  K2j  K'ubK(j  )��}�(h�jP  j  ]�j  K2j  K(ubK)j  )��}�(h�jP  j  ]�j  K2j  K)ubK*j  )��}�(h�jP  j  ]�j  K2j  K*ubK+j  )��}�(h�jP  j  ]�j  K2j  K+ubK,j  )��}�(h�jP  j  ]�j  K2j  K,ubK-j  )��}�(h�jP  j  ]�j  K2j  K-ubK.j  )��}�(h�jP  j  ]�j  K2j  K.ubK/j  )��}�(h�jP  j  ]�j  K2j  K/ubK0j  )��}�(h�jP  j  ]�j  K2j  K0ubK1j  )��}�(h�jP  j  ]�j  K2j  K1ubK2j  )��}�(h�jP  j  ]�j  K2j  K2ubK3j  )��}�(h�jP  j  ]�j  K2j  K3ubK4j  )��}�(h�jP  j  ]�j  K2j  K4ubK5j  )��}�(h�jP  j  ]�j  K2j  K5ubK6j  )��}�(h�jP  j  ]�j  K2j  K6ubK7j  )��}�(h�jP  j  ]�j  K2j  K7ubK8j  )��}�(h�jP  j  ]�j  K2j  K8ubK9j  )��}�(h�jP  j  ]�j  K2j  K9ubK:j  )��}�(h�jP  j  ]�j  K2j  K:ubK;j  )��}�(h�jP  j  ]�j  K2j  K;ubuK3}�(K j  )��}�(h�jP  j  ]�j  K3j  K ubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubK	j  )��}�(h�jP  j  ]�j  K3j  K	ubK
j  )��}�(h�jP  j  ]�j  K3j  K
ubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubKj  )��}�(h�jP  j  ]�j  K3j  KubK j  )��}�(h�jP  j  ]�j  K3j  K ubK!j  )��}�(h�jP  j  ]�j  K3j  K!ubK"j  )��}�(h�jP  j  ]�j  K3j  K"ubK#j  )��}�(h�jP  j  ]�j  K3j  K#ubK$j  )��}�(h�jP  j  ]�j  K3j  K$ubK%j  )��}�(h�jP  j  ]�j  K3j  K%ubK&j  )��}�(h�jP  j  ]�j  K3j  K&ubK'j  )��}�(h�jP  j  ]�j  K3j  K'ubK(j  )��}�(h�jP  j  ]�j  K3j  K(ubK)j  )��}�(h�jP  j  ]�j  K3j  K)ubK*j  )��}�(h�jP  j  ]�j  K3j  K*ubK+j  )��}�(h�jP  j  ]�j  K3j  K+ubK,j  )��}�(h�jP  j  ]�j  K3j  K,ubK-j  )��}�(h�jP  j  ]�j  K3j  K-ubK.j  )��}�(h�jP  j  ]�j  K3j  K.ubK/j  )��}�(h�jP  j  ]�j  K3j  K/ubK0j  )��}�(h�jP  j  ]�j  K3j  K0ubK1j  )��}�(h�jP  j  ]�j  K3j  K1ubK2j  )��}�(h�jP  j  ]�j  K3j  K2ubK3j  )��}�(h�jP  j  ]�j  K3j  K3ubK4j  )��}�(h�jP  j  ]�j  K3j  K4ubK5j  )��}�(h�jP  j  ]�j  K3j  K5ubK6j  )��}�(h�jP  j  ]�j  K3j  K6ubK7j  )��}�(h�jP  j  ]�j  K3j  K7ubK8j  )��}�(h�jP  j  ]�j  K3j  K8ubK9j  )��}�(h�jP  j  ]�j  K3j  K9ubK:j  )��}�(h�jP  j  ]�j  K3j  K:ubK;j  )��}�(h�jP  j  ]�j  K3j  K;ubuK4}�(K j  )��}�(h�jP  j  ]�j  K4j  K ubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubK	j  )��}�(h�jP  j  ]�j  K4j  K	ubK
j  )��}�(h�jP  j  ]�j  K4j  K
ubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubKj  )��}�(h�jP  j  ]�j  K4j  KubK j  )��}�(h�jP  j  ]�j  K4j  K ubK!j  )��}�(h�jP  j  ]�j  K4j  K!ubK"j  )��}�(h�jP  j  ]�j  K4j  K"ubK#j  )��}�(h�jP  j  ]�j  K4j  K#ubK$j  )��}�(h�jP  j  ]�j  K4j  K$ubK%j  )��}�(h�jP  j  ]�j  K4j  K%ubK&j  )��}�(h�jP  j  ]�j  K4j  K&ubK'j  )��}�(h�jP  j  ]�j  K4j  K'ubK(j  )��}�(h�jP  j  ]�j  K4j  K(ubK)j  )��}�(h�jP  j  ]�j  K4j  K)ubK*j  )��}�(h�jP  j  ]�j  K4j  K*ubK+j  )��}�(h�jP  j  ]�j  K4j  K+ubK,j  )��}�(h�jP  j  ]�j  K4j  K,ubK-j  )��}�(h�jP  j  ]�j  K4j  K-ubK.j  )��}�(h�jP  j  ]�j  K4j  K.ubK/j  )��}�(h�jP  j  ]�j  K4j  K/ubK0j  )��}�(h�jP  j  ]�j  K4j  K0ubK1j  )��}�(h�jP  j  ]�j  K4j  K1ubK2j  )��}�(h�jP  j  ]�j  K4j  K2ubK3j  )��}�(h�jP  j  ]�j  K4j  K3ubK4j  )��}�(h�jP  j  ]�j  K4j  K4ubK5j  )��}�(h�jP  j  ]�j  K4j  K5ubK6j  )��}�(h�jP  j  ]�j  K4j  K6ubK7j  )��}�(h�jP  j  ]�j  K4j  K7ubK8j  )��}�(h�jP  j  ]�j  K4j  K8ubK9j  )��}�(h�jP  j  ]�j  K4j  K9ubK:j  )��}�(h�jP  j  ]�j  K4j  K:ubK;j  )��}�(h�jP  j  ]�j  K4j  K;ubuK5}�(K j  )��}�(h�jP  j  ]�j  K5j  K ubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubK	j  )��}�(h�jP  j  ]�j  K5j  K	ubK
j  )��}�(h�jP  j  ]�j  K5j  K
ubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubKj  )��}�(h�jP  j  ]�j  K5j  KubK j  )��}�(h�jP  j  ]�j  K5j  K ubK!j  )��}�(h�jP  j  ]�j  K5j  K!ubK"j  )��}�(h�jP  j  ]�j  K5j  K"ubK#j  )��}�(h�jP  j  ]�j  K5j  K#ubK$j  )��}�(h�jP  j  ]�j  K5j  K$ubK%j  )��}�(h�jP  j  ]�j  K5j  K%ubK&j  )��}�(h�jP  j  ]�j  K5j  K&ubK'j  )��}�(h�jP  j  ]�j  K5j  K'ubK(j  )��}�(h�jP  j  ]�j  K5j  K(ubK)j  )��}�(h�jP  j  ]�j  K5j  K)ubK*j  )��}�(h�jP  j  ]�j  K5j  K*ubK+j  )��}�(h�jP  j  ]�j  K5j  K+ubK,j  )��}�(h�jP  j  ]�j  K5j  K,ubK-j  )��}�(h�jP  j  ]�j  K5j  K-ubK.j  )��}�(h�jP  j  ]�j  K5j  K.ubK/j  )��}�(h�jP  j  ]�j  K5j  K/ubK0j  )��}�(h�jP  j  ]�j  K5j  K0ubK1j  )��}�(h�jP  j  ]�j  K5j  K1ubK2j  )��}�(h�jP  j  ]�j  K5j  K2ubK3j  )��}�(h�jP  j  ]�j  K5j  K3ubK4j  )��}�(h�jP  j  ]�j  K5j  K4ubK5j  )��}�(h�jP  j  ]�j  K5j  K5ubK6j  )��}�(h�jP  j  ]�j  K5j  K6ubK7j  )��}�(h�jP  j  ]�j  K5j  K7ubK8j  )��}�(h�jP  j  ]�j  K5j  K8ubK9j  )��}�(h�jP  j  ]�j  K5j  K9ubK:j  )��}�(h�jP  j  ]�j  K5j  K:ubK;j  )��}�(h�jP  j  ]�j  K5j  K;ubuK6}�(K j  )��}�(h�jP  j  ]�j  K6j  K ubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubK	j  )��}�(h�jP  j  ]�j  K6j  K	ubK
j  )��}�(h�jP  j  ]�j  K6j  K
ubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubKj  )��}�(h�jP  j  ]�j  K6j  KubK j  )��}�(h�jP  j  ]�j  K6j  K ubK!j  )��}�(h�jP  j  ]�j  K6j  K!ubK"j  )��}�(h�jP  j  ]�j  K6j  K"ubK#j  )��}�(h�jP  j  ]�j  K6j  K#ubK$j  )��}�(h�jP  j  ]�j  K6j  K$ubK%j  )��}�(h�jP  j  ]�j  K6j  K%ubK&j  )��}�(h�jP  j  ]�j  K6j  K&ubK'j  )��}�(h�jP  j  ]�j  K6j  K'ubK(j  )��}�(h�jP  j  ]�j  K6j  K(ubK)j  )��}�(h�jP  j  ]�j  K6j  K)ubK*j  )��}�(h�jP  j  ]�j  K6j  K*ubK+j  )��}�(h�jP  j  ]�j  K6j  K+ubK,j  )��}�(h�jP  j  ]�j  K6j  K,ubK-j  )��}�(h�jP  j  ]�j  K6j  K-ubK.j  )��}�(h�jP  j  ]�j  K6j  K.ubK/j  )��}�(h�jP  j  ]�j  K6j  K/ubK0j  )��}�(h�jP  j  ]�j  K6j  K0ubK1j  )��}�(h�jP  j  ]�j  K6j  K1ubK2j  )��}�(h�jP  j  ]�j  K6j  K2ubK3j  )��}�(h�jP  j  ]�j  K6j  K3ubK4j  )��}�(h�jP  j  ]�j  K6j  K4ubK5j  )��}�(h�jP  j  ]�j  K6j  K5ubK6j  )��}�(h�jP  j  ]�j  K6j  K6ubK7j  )��}�(h�jP  j  ]�j  K6j  K7ubK8j  )��}�(h�jP  j  ]�j  K6j  K8ubK9j  )��}�(h�jP  j  ]�j  K6j  K9ubK:j  )��}�(h�jP  j  ]�j  K6j  K:ubK;j  )��}�(h�jP  j  ]�j  K6j  K;ubuK7}�(K j  )��}�(h�jP  j  ]�j  K7j  K ubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubK	j  )��}�(h�jP  j  ]�j  K7j  K	ubK
j  )��}�(h�jP  j  ]�j  K7j  K
ubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubKj  )��}�(h�jP  j  ]�j  K7j  KubK j  )��}�(h�jP  j  ]�j  K7j  K ubK!j  )��}�(h�jP  j  ]�j  K7j  K!ubK"j  )��}�(h�jP  j  ]�j  K7j  K"ubK#j  )��}�(h�jP  j  ]�j  K7j  K#ubK$j  )��}�(h�jP  j  ]�j  K7j  K$ubK%j  )��}�(h�jP  j  ]�j  K7j  K%ubK&j  )��}�(h�jP  j  ]�j  K7j  K&ubK'j  )��}�(h�jP  j  ]�j  K7j  K'ubK(j  )��}�(h�jP  j  ]�j  K7j  K(ubK)j  )��}�(h�jP  j  ]�j  K7j  K)ubK*j  )��}�(h�jP  j  ]�j  K7j  K*ubK+j  )��}�(h�jP  j  ]�j  K7j  K+ubK,j  )��}�(h�jP  j  ]�j  K7j  K,ubK-j  )��}�(h�jP  j  ]�j  K7j  K-ubK.j  )��}�(h�jP  j  ]�j  K7j  K.ubK/j  )��}�(h�jP  j  ]�j  K7j  K/ubK0j  )��}�(h�jP  j  ]�j  K7j  K0ubK1j  )��}�(h�jP  j  ]�j  K7j  K1ubK2j  )��}�(h�jP  j  ]�j  K7j  K2ubK3j  )��}�(h�jP  j  ]�j  K7j  K3ubK4j  )��}�(h�jP  j  ]�j  K7j  K4ubK5j  )��}�(h�jP  j  ]�j  K7j  K5ubK6j  )��}�(h�jP  j  ]�j  K7j  K6ubK7j  )��}�(h�jP  j  ]�j  K7j  K7ubK8j  )��}�(h�jP  j  ]�j  K7j  K8ubK9j  )��}�(h�jP  j  ]�j  K7j  K9ubK:j  )��}�(h�jP  j  ]�j  K7j  K:ubK;j  )��}�(h�jP  j  ]�j  K7j  K;ubuK8}�(K j  )��}�(h�jP  j  ]�j  K8j  K ubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubK	j  )��}�(h�jP  j  ]�j  K8j  K	ubK
j  )��}�(h�jP  j  ]�j  K8j  K
ubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubKj  )��}�(h�jP  j  ]�j  K8j  KubK j  )��}�(h�jP  j  ]�j  K8j  K ubK!j  )��}�(h�jP  j  ]�j  K8j  K!ubK"j  )��}�(h�jP  j  ]�j  K8j  K"ubK#j  )��}�(h�jP  j  ]�j  K8j  K#ubK$j  )��}�(h�jP  j  ]�j  K8j  K$ubK%j  )��}�(h�jP  j  ]�j  K8j  K%ubK&j  )��}�(h�jP  j  ]�j  K8j  K&ubK'j  )��}�(h�jP  j  ]�j  K8j  K'ubK(j  )��}�(h�jP  j  ]�j  K8j  K(ubK)j  )��}�(h�jP  j  ]�j  K8j  K)ubK*j  )��}�(h�jP  j  ]�j  K8j  K*ubK+j  )��}�(h�jP  j  ]�j  K8j  K+ubK,j  )��}�(h�jP  j  ]�j  K8j  K,ubK-j  )��}�(h�jP  j  ]�j  K8j  K-ubK.j  )��}�(h�jP  j  ]�j  K8j  K.ubK/j  )��}�(h�jP  j  ]�j  K8j  K/ubK0j  )��}�(h�jP  j  ]�j  K8j  K0ubK1j  )��}�(h�jP  j  ]�j  K8j  K1ubK2j  )��}�(h�jP  j  ]�j  K8j  K2ubK3j  )��}�(h�jP  j  ]�j  K8j  K3ubK4j  )��}�(h�jP  j  ]�j  K8j  K4ubK5j  )��}�(h�jP  j  ]�j  K8j  K5ubK6j  )��}�(h�jP  j  ]�j  K8j  K6ubK7j  )��}�(h�jP  j  ]�j  K8j  K7ubK8j  )��}�(h�jP  j  ]�j  K8j  K8ubK9j  )��}�(h�jP  j  ]�j  K8j  K9ubK:j  )��}�(h�jP  j  ]�j  K8j  K:ubK;j  )��}�(h�jP  j  ]�j  K8j  K;ubuK9}�(K j  )��}�(h�jP  j  ]�j  K9j  K ubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubK	j  )��}�(h�jP  j  ]�j  K9j  K	ubK
j  )��}�(h�jP  j  ]�j  K9j  K
ubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubKj  )��}�(h�jP  j  ]�j  K9j  KubK j  )��}�(h�jP  j  ]�j  K9j  K ubK!j  )��}�(h�jP  j  ]�j  K9j  K!ubK"j  )��}�(h�jP  j  ]�j  K9j  K"ubK#j  )��}�(h�jP  j  ]�j  K9j  K#ubK$j  )��}�(h�jP  j  ]�j  K9j  K$ubK%j  )��}�(h�jP  j  ]�j  K9j  K%ubK&j  )��}�(h�jP  j  ]�j  K9j  K&ubK'j  )��}�(h�jP  j  ]�j  K9j  K'ubK(j  )��}�(h�jP  j  ]�j  K9j  K(ubK)j  )��}�(h�jP  j  ]�j  K9j  K)ubK*j  )��}�(h�jP  j  ]�j  K9j  K*ubK+j  )��}�(h�jP  j  ]�j  K9j  K+ubK,j  )��}�(h�jP  j  ]�j  K9j  K,ubK-j  )��}�(h�jP  j  ]�j  K9j  K-ubK.j  )��}�(h�jP  j  ]�j  K9j  K.ubK/j  )��}�(h�jP  j  ]�j  K9j  K/ubK0j  )��}�(h�jP  j  ]�j  K9j  K0ubK1j  )��}�(h�jP  j  ]�j  K9j  K1ubK2j  )��}�(h�jP  j  ]�j  K9j  K2ubK3j  )��}�(h�jP  j  ]�j  K9j  K3ubK4j  )��}�(h�jP  j  ]�j  K9j  K4ubK5j  )��}�(h�jP  j  ]�j  K9j  K5ubK6j  )��}�(h�jP  j  ]�j  K9j  K6ubK7j  )��}�(h�jP  j  ]�j  K9j  K7ubK8j  )��}�(h�jP  j  ]�j  K9j  K8ubK9j  )��}�(h�jP  j  ]�j  K9j  K9ubK:j  )��}�(h�jP  j  ]�j  K9j  K:ubK;j  )��}�(h�jP  j  ]�j  K9j  K;ubuK:}�(K j  )��}�(h�jP  j  ]�j  K:j  K ubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubK	j  )��}�(h�jP  j  ]�j  K:j  K	ubK
j  )��}�(h�jP  j  ]�j  K:j  K
ubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubKj  )��}�(h�jP  j  ]�j  K:j  KubK j  )��}�(h�jP  j  ]�j  K:j  K ubK!j  )��}�(h�jP  j  ]�j  K:j  K!ubK"j  )��}�(h�jP  j  ]�j  K:j  K"ubK#j  )��}�(h�jP  j  ]�j  K:j  K#ubK$j  )��}�(h�jP  j  ]�j  K:j  K$ubK%j  )��}�(h�jP  j  ]�j  K:j  K%ubK&j  )��}�(h�jP  j  ]�j  K:j  K&ubK'j  )��}�(h�jP  j  ]�j  K:j  K'ubK(j  )��}�(h�jP  j  ]�j  K:j  K(ubK)j  )��}�(h�jP  j  ]�j  K:j  K)ubK*j  )��}�(h�jP  j  ]�j  K:j  K*ubK+j  )��}�(h�jP  j  ]�j  K:j  K+ubK,j  )��}�(h�jP  j  ]�j  K:j  K,ubK-j  )��}�(h�jP  j  ]�j  K:j  K-ubK.j  )��}�(h�jP  j  ]�j  K:j  K.ubK/j  )��}�(h�jP  j  ]�j  K:j  K/ubK0j  )��}�(h�jP  j  ]�j  K:j  K0ubK1j  )��}�(h�jP  j  ]�j  K:j  K1ubK2j  )��}�(h�jP  j  ]�j  K:j  K2ubK3j  )��}�(h�jP  j  ]�j  K:j  K3ubK4j  )��}�(h�jP  j  ]�j  K:j  K4ubK5j  )��}�(h�jP  j  ]�j  K:j  K5ubK6j  )��}�(h�jP  j  ]�j  K:j  K6ubK7j  )��}�(h�jP  j  ]�j  K:j  K7ubK8j  )��}�(h�jP  j  ]�j  K:j  K8ubK9j  )��}�(h�jP  j  ]�j  K:j  K9ubK:j  )��}�(h�jP  j  ]�j  K:j  K:ubK;j  )��}�(h�jP  j  ]�j  K:j  K;ubuK;}�(K j  )��}�(h�jP  j  ]�j  K;j  K ubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubK	j  )��}�(h�jP  j  ]�j  K;j  K	ubK
j  )��}�(h�jP  j  ]�j  K;j  K
ubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubKj  )��}�(h�jP  j  ]�j  K;j  KubK j  )��}�(h�jP  j  ]�j  K;j  K ubK!j  )��}�(h�jP  j  ]�j  K;j  K!ubK"j  )��}�(h�jP  j  ]�j  K;j  K"ubK#j  )��}�(h�jP  j  ]�j  K;j  K#ubK$j  )��}�(h�jP  j  ]�j  K;j  K$ubK%j  )��}�(h�jP  j  ]�j  K;j  K%ubK&j  )��}�(h�jP  j  ]�j  K;j  K&ubK'j  )��}�(h�jP  j  ]�j  K;j  K'ubK(j  )��}�(h�jP  j  ]�j  K;j  K(ubK)j  )��}�(h�jP  j  ]�j  K;j  K)ubK*j  )��}�(h�jP  j  ]�j  K;j  K*ubK+j  )��}�(h�jP  j  ]�j  K;j  K+ubK,j  )��}�(h�jP  j  ]�j  K;j  K,ubK-j  )��}�(h�jP  j  ]�j  K;j  K-ubK.j  )��}�(h�jP  j  ]�j  K;j  K.ubK/j  )��}�(h�jP  j  ]�j  K;j  K/ubK0j  )��}�(h�jP  j  ]�j  K;j  K0ubK1j  )��}�(h�jP  j  ]�j  K;j  K1ubK2j  )��}�(h�jP  j  ]�j  K;j  K2ubK3j  )��}�(h�jP  j  ]�j  K;j  K3ubK4j  )��}�(h�jP  j  ]�j  K;j  K4ubK5j  )��}�(h�jP  j  ]�j  K;j  K5ubK6j  )��}�(h�jP  j  ]�j  K;j  K6ubK7j  )��}�(h�jP  j  ]�j  K;j  K7ubK8j  )��}�(h�jP  j  ]�j  K;j  K8ubK9j  )��}�(h�jP  j  ]�j  K;j  K9ubK:j  )��}�(h�jP  j  ]�j  K;j  K:ubK;j  )��}�(h�jP  j  ]�j  K;j  K;ubuujcN  jdN  jeN  ]�(]�(K'K'e]�(K&K&e]�(K'K)e]�(K&K*e]�(K'K'e]�(K&K&e]�(K'K)e]�(K&K*e]�(K'K'e]�(K&K&e]�(K'K)e]�(K&K*e]�(K'K'e]�(K&K&e]�(K'K)e]�(K'K*e]�(K'K'e]�(K'K&e]�(K&K%e]�(K'K)e]�(K'K*e]�(K'K'e]�(K'K&e]�(K&K%e]�(K'K)e]�(K'K*e]�(K'K'e]�(K'K&e]�(K&K%e]�(K(K)e]�(K'K*e]�(K(K'e]�(K'K&e]�(K'K%e]�(K(K)e]�(K'K*e]�(K(K'e]�(K'K&e]�(K'K%e]�(K(K)e]�(K'K*e]�(K(K'e]�(K'K&e]�(K'K%e]�(K(K)e]�(K(K*e]�(K(K'e]�(K(K&e]�(K'K%e]�(K(K)e]�(K(K*e]�(K(K'e]�(K(K&e]�(K(K%e]�(K(K$e]�(K(K)e]�(K(K*e]�(K(K'e]�(K(K&e]�(K(K%e]�(K(K$e]�(K(K)e]�(K(K*e]�(K(K'e]�(K(K&e]�(K(K%e]�(K(K$e]�(K(K)e]�(K(K*e]�(K(K'e]�(K(K&e]�(K)K%e]�(K)K$e]�(K)K#e]�(K(K)e]�(K(K*e]�(K(K'e]�(K)K&e]�(K)K%e]�(K)K$e]�(K)K#e]�(K(K)e]�(K(K*e]�(K(K'e]�(K)K&e]�(K)K%e]�(K)K$e]�(K*K#e]�(K(K)e]�(K)K*e]�(K(K'e]�(K)K&e]�(K)K%e]�(K*K$e]�(K*K#e]�(K(K)e]�(K)K*e]�(K)K'e]�(K)K&e]�(K*K%e]�(K*K$e]�(K+K#e]�(K(K)e]�(K)K*e]�(K)K'e]�(K)K&e]�(K*K%e]�(K*K$e]�(K+K#e]�(K)K)e]�(K)K*e]�(K)K'e]�(K)K&e]�(K*K%e]�(K+K$e]�(K+K#e]�(K)K)e]�(K)K*e]�(K)K'e]�(K*K&e]�(K*K%e]�(K+K$e]�(K,K#e]�(K-K"e]�(K)K)e]�(K)K*e]�(K)K'e]�(K*K&e]�(K+K%e]�(K+K$e]�(K,K#e]�(K-K"e]�(K)K)e]�(K*K*e]�(K)K'e]�(K*K&e]�(K+K%e]�(K,K$e]�(K-K#e]�(K)K)e]�(K*K*e]�(K)K'e]�(K*K&e]�(K+K%e]�(K,K$e]�(K-K#e]�(K)K)e]�(K*K*e]�(K'K'e]�(K&K&e]�(K)K'e]�(K*K&e]�(K+K%e]�(K,K$e]�(K-K#e]�(K'K'e]�(K&K&e]�(K)K'e]�(K*K&e]�(K+K%e]�(K,K$e]�(K-K#e]�(K'K'e]�(K&K&e]�(K)K'e]�(K*K&e]�(K+K&e]�(K,K%e]�(K-K$e]�(K.K#e]�(K'K'e]�(K&K&e]�(K)K'e]�(K*K'e]�(K+K&e]�(K,K%e]�(K-K$e]�(K.K$e]�(K/K#e]�(K'K'e]�(K&K'e]�(K)K'e]�(K*K'e]�(K+K&e]�(K,K%e]�(K-K%e]�(K.K$e]�(K/K#e]�(K'K'e]�(K&K'e]�(K)K'e]�(K*K'e]�(K+K&e]�(K,K&e]�(K-K%e]�(K.K%e]�(K/K$e]�(K0K#e]�(K'K'e]�(K&K'e]�(K)K(e]�(K*K'e]�(K+K'e]�(K,K&e]�(K-K&e]�(K.K%e]�(K/K%e]�(K0K$e]�(K'K(e]�(K&K'e]�(K)K(e]�(K*K'e]�(K+K'e]�(K,K&e]�(K-K&e]�(K.K&e]�(K/K%e]�(K0K%e]�(K'K(e]�(K&K'e]�(K)K(e]�(K*K'e]�(K+K'e]�(K,K'e]�(K-K&e]�(K.K&e]�(K/K&e]�(K0K%e]�(K'K(e]�(K&K'e]�(K)K(e]�(K*K(e]�(K+K'e]�(K,K'e]�(K-K'e]�(K.K'e]�(K/K&e]�(K0K&e]�(K'K(e]�(K&K(e]�(K)K(e]�(K*K(e]�(K+K(e]�(K,K'e]�(K-K'e]�(K.K'e]�(K/K'e]�(K0K'e]�(K'K(e]�(K&K(e]�(K)K(e]�(K*K(e]�(K+K(e]�(K,K(e]�(K-K(e]�(K.K(e]�(K/K'e]�(K0K'e]�(K'K(e]�(K&K(e]�(K)K(e]�(K*K(e]�(K+K(e]�(K,K(e]�(K-K(e]�(K.K(e]�(K/K(e]�(K0K(e]�(K'K(e]�(K&K(e]�(K)K(e]�(K*K(e]�(K+K(e]�(K,K(e]�(K-K(e]�(K.K(e]�(K/K)e]�(K0K)e]�(K'K(e]�(K&K(e]�(K)K(e]�(K*K(e]�(K+K(e]�(K,K)e]�(K-K)e]�(K.K)e]�(K/K)e]�(K0K)e]�(K'K(e]�(K&K)e]�(K)K(e]�(K*K(e]�(K+K)e]�(K,K)e]�(K-K)e]�(K.K)e]�(K/K*e]�(K'K(e]�(K&K)e]�(K)K(e]�(K*K)e]�(K+K)e]�(K,K)e]�(K-K*e]�(K'K(e]�(K&K)e]�(K)K(e]�(K*K)e]�(K+K)e]�(K,K*e]�(K'K)e]�(K&K)e]�(K)K(e]�(K*K)e]�(K+K)e]�(K,K*e]�(K'K)e]�(K&K)e]�(K)K)e]�(K*K)e]�(K+K*e]�(K'K)e]�(K&K)e]�(K)K)e]�(K*K)e]�(K+K*e]�(K'K)e]�(K&K*e]�(K)K)e]�(K*K)e]�(K+K*e]�(K'K)e]�(K&K*e]�(K)K)e]�(K*K*e]�(K'K)e]�(K&K*e]�(K)K)e]�(K*K*e]�(K'K)e]�(K&K*e]�(K)K)e]�(K*K*e]�(K(K(e]�(K(K)eeh[jYP  j	O  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNG�`�     G�`�     G�`�     G�`�     NNNNNNNNNNNG�b�     G�c      G�cP     G�c�     G�c�     G�c�     G�d     G�d@     G�dp     G�d�     G�d�     G�e      G�d�     G�d�     G�dp     G�d�     G�d�     G�e      K NNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�`�     G�`�     G�`�     G�`P     G�`�     NNNNNNNNNNNG�b�     NNNNNNNNNNG�d�     G�d�     G�dp     G�d@     G�dp     G�d�     G�d�     G�e      NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`�     G�`�     G�`P     G�`      G�`P     NNNNNNNNNNNG�b�     NNNNNNNNNNG�d�     G�dp     G�d@     G�d     G�d@     G�dp     G�d�     G�d�     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`�     G�`P     G�`      G�_�     G�`      NNNNNNNNNNNG�b`     NNNNNNNNNNG�dp     G�d@     G�d     G�c�     G�d     G�d@     G�dp     G�d�     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`P     G�`      G�_�     G�_�     G�_�     NNNNNNNNNNNG�b0     NNNNNNNNNNNG�d     G�c�     G�c�     G�c�     G�d     G�d@     G�dp     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`P     G�`      G�_�     G�_�     G�_      G�_�     G�_�     G�`      G�`P     G�`�     G�`�     G�`�     G�a     G�a@     G�ap     G�a�     G�a�     G�b      NNNNNNNNNNNNG�c�     G�c�     G�c�     G�c�     G�d     G�d@     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`      G�_�     G�_�     G�_      G�^�     G�_      NNNNNNNNNNNNNNNNNNNNNNNNNG�cP     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�_�     G�_�     G�_      G�^�     G�^`     G�^�     NNNNNNNNNNNNNNNNNNNNNNNNNG�c      NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�_�     G�_      G�^�     G�^`     G�^      G�^`     NNNNNNNNNNNNNNNNNNNNNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�]�     NNNNNNNNNNNNNNNNNNNNNNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�]@     NNNNNNNNNNNNNNNNNNNNNNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�\�     NNNNNNNNNNNNNNNNNNNNNNNNNNG�b`     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�\�     NNNNNNNNNNNNNNNNNNNNNNNNNNG�b0     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�\      NNNNNNNNNNNNNNNNNNNNNNNNNNG�b      NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�[�     G�[`     G�[      G�Z�     NNNNNNNNNNNNNNNNNNNNNNNG�a�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�Z@     NNNNNNNNNNNNNNNNNNNNNNNG�a�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�Y�     NNNNNNNNNNNNNNNNNNNNNNNG�ap     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�Y�     NNNNNNNNNNNNNNNNNNNNNNNG�a@     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�Y      NNNNNNNNNNNNNNNNNNNNNNNG�a     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�X�     NNNNNNNNNNNNNNNNNNNNNNNG�`�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�X`     NNNNNNNNNNNNNG�]�     G�^      G�^`     G�^�     G�_      G�_�     G�_�     G�`      G�`P     G�`�     G�`�     G�`�     G�a     G�a@     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�X      NNNNNNNNNNNNNG�]@     NNNNNNG�`P     G�`�     G�`�     G�`�     G�a     G�a@     G�ap     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�V�     G�W@     G�W�     G�X      G�X`     G�X�     NNNNNNNNNNG�\�     NNNNNNG�`�     G�`�     G�`�     G�a     G�a@     G�ap     G�a�     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�V�     G�V�     G�W@     G�W�     G�X      G�X`     NNNNNNNNNNG�\�     NNNNNNG�`�     G�`�     G�a     G�a@     G�ap     G�a�     G�a�     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�V      G�V�     G�V�     G�W@     G�W�     G�X      NNNNNNNNNNG�\      NNNNNNG�`�     G�a     G�a@     G�ap     G�a�     G�a�     G�b      NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�U�     G�V      G�V�     G�V�     G�W@     G�W�     G�X      G�X`     G�X�     G�Y      G�Y�     G�Y�     G�Z@     G�Z�     G�[      G�[`     G�[�     NNNNNNG�a     G�a@     G�ap     G�a�     G�a�     G�b      G�b0     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�U`     G�U�     G�V      G�V�     G�V�     G�W@     NNNNNNNNNNNNNNNNNG�a@     G�ap     G�a�     G�a�     G�b      G�b0     G�b`     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�U      G�U`     G�U�     G�V      G�V�     G�V�     NNNNNNNNNNNNNNNNNG�ap     G�a�     G�a�     G�b      G�b0     G�b`     G�b�     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�T�     G�U      G�U`     G�U�     G�V      G�V�     NNNNNNNNNNNNNNNNNG�a�     G�a�     G�b      G�b0     G�b`     G�b�     G�b�     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�T@     G�T�     G�U      G�U`     G�U�     G�V      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�S�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�S�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�S      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�R�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�R`     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNG�P�     G�Q@     G�Q�     G�R      NNNNNNNNNNNNNNNNNNNNNNNNNNN�      NNNG�      G�      G��      G�      NNNNNNNNNNNNNNNNNNe]�(NNNNG�P�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�      G�      G��      G�       G��      NNNNNNNNNNNNNNNNNNe]�(NNNNG�P      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�      G�      G�      G�      G��      G�      NNNNNNNNNNNNNNNNNNe]�(NNNNG�O�     G�N�     G�N      G�M@     G�L�     NNNNNNNNNNNNNNNNNNNNNNNNNNNG�"      G�      G�      G�      G�      G�      NNNNNNNNNNNNNNNNNNe]�(NNNNG�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     NNNNNNNNNNNNNNNNG�%      G�"      G�      G�      G�      G�      NNNNNNNNNNNNNNNNNNe]�(NNNNG�O�     G�N�     G�N      G�M@     G�L�     NNNNNNNNNNG�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�(      G�%      G�"      G�      G�      G�      NNNNNNNNNNNNNNNNNNe]�(NNNNG�P      G�O�     G�N�     G�N      G�M@     NNNNNNNNNNNNNNNNNNNNNNNNNNNG�+      G�(      G�%      G�"      G�      G�"      NNNNNNNNNNNNNNNNNNe]�(NNNNG�P�     G�P      G�O�     G�N�     G�N      NNNNNNNNNNNNNNNNNNNNNNNNNNNG�.      G�+      G�(      G�%      G�"      G�%      NNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�0�     G�.      G�+      G�(      G�%      G�(      NNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej[O  ]�(j�  jo  j  ej]O  j^O  j_O  ]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K eej�O  ]�(]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  jl  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jM  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  hUj�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jM  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jM  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  jA  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jl  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jM  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  hUj�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jl  j�O  j�O  j�O  j~  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j  jM  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  jM  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  e]�(j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  j�O  eejP  jP  �	thePlayer�h�consumeList�]�(hQh�h�h�hre�	tilesSeen�]��
stairsDown�]�(K(K)e�djikstra_Stairs_Up�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKKKKNNNNNNNNNNNKKKKKKKKKKKKK K!K"K#K$K%K&NNNNNNNNNNNNNNNNNNNNNNe]�(NNNKKKKKNNNNNNNNNNNKNNNNNNNNNNK K!K"K#K$K%K&K'NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNKNNNNNNNNNNK!K"K#K$K%K&K'K(NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKK KNNNNNNNNNNNKNNNNNNNNNNK"K#K$K%K&K'K(K)NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNKNNNNNNNNNNNK$K%K&K'K(K)K*NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKKKKKKK	K
KKKKKNNNNNNNNNNNNK&K'K(K)K*K+NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNK(NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNK)NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK	KKKKKNNNNNNNNNNNNNNNNNNNNNNNNNK*NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK+NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK,NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK-NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK	NNNNNNNNNNNNNNNNNNNNNNNNNNK.NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK
NNNNNNNNNNNNNNNNNNNNNNNNNNK/NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKKKKNNNNNNNNNNNNNNNNNNNNNNNK0NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK5NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNK,K-K.K/K0K1K2K3K4K5K6K7K8K9NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNK+NNNNNNK4K5K6K7K8K9K:NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNK*NNNNNNK5K6K7K8K9K:K;NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNK)NNNNNNK6K7K8K9K:K;K<NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNK(NNNNNNK7K8K9K:K;K<K=NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKKKKK K!K"K#K$K%K&K'NNNNNNK8K9K:K;K<K=K>NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNK9K:K;K<K=K>K?NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNK:K;K<K=K>K?K@NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNK;K<K=K>K?K@KANNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKK NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK!NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK"NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK#NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK$NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNK(K'K&K%NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKTKUKVKWNNNNNNNNNNNNNNNNNNe]�(NNNNK)NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKRKSKTKUKVNNNNNNNNNNNNNNNNNNe]�(NNNNK*NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKPKQKRKSKTKUNNNNNNNNNNNNNNNNNNe]�(NNNNK+K,K-K.K/NNNNNNNNNNNNNNNNNNNNNNNNNNNKOKPKQKRKSKTNNNNNNNNNNNNNNNNNNe]�(NNNNK,K-K.K/K0K1K2K3K4K5K6K7K8K9K:K;NNNNNNNNNNNNNNNNKNKOKPKQKRKSNNNNNNNNNNNNNNNNNNe]�(NNNNK-K.K/K0K1NNNNNNNNNNK<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQKRNNNNNNNNNNNNNNNNNNe]�(NNNNK.K/K0K1K2NNNNNNNNNNNNNNNNNNNNNNNNNNNKNKOKPKQKRKSNNNNNNNNNNNNNNNNNNe]�(NNNNK/K0K1K2K3NNNNNNNNNNNNNNNNNNNNNNNNNNNKOKPKQKRKSKTNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKPKQKRKSKTKUNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�	gameState��__main__��Game���)��}�(�loadRequest���console��tdl��Console���)��KYK*]�(K K K K ��K K K ����KKK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KLK�K�K���K K K ����KEK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KRK�K�K���K K K ����KPK�K�K���K K K ����KAK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KWK�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KSK�K�K���K K K ����KSK�K�K���K K K ����KZK�K�K���K K K ����KKK�K�K���K K K ����K-K�K�K���K K K ����KKK�K�K���K K K ����KZK�K�K���K K K ����KKK�K�K���K K K ����KZK�K�K���K K K ����KZK�K�K���K K K ����KZK�K�K���K K K ����KZK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KxK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KaK�K�K���K K K ����KoK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KoK�K�K���K K K ����KyK�K�K���K K K ����K-K�K�K���K K K ����KyK�K�K���K K K ����KoK�K�K���K K K ����KyK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����KFK�K�K���K K K ����K K K K ��K K K ����KvK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KnK�K�K���K K K ����KwK�K�K���K K K ����KmK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KmK�K�K���K K K ����KlK�K�K���K K K ����K-K�K�K���K K K ����KlK�K�K���K K K ����KmK�K�K���K K K ����KlK�K�K���K K K ����KmK�K�K���K K K ����KmK�K�K���K K K ����KmK�K�K���K K K ����KmK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KbK�K�K���K K K ����KeK�K�K���K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KbK�K�K���K K K ����KeK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KwK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KiK�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����KiK�K�K���K K K ����K K�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K3K�K�K���K K K ����K K K K ��K K K ����KhK�K�K���K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K:K�K�K���K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����KeK�K�K���K K K ����KpK�K�K���K K K ����K-K�K�K���K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KPK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K6K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����KiK�K�K���K K K ����K-K�K�K���K K K ����KtK�K�K���K K K ����K K�K�K���K K K ����KtK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KcK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K1K�K�K���K K K ����K4K�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K7K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����KcK�K�K���K K K ����K-K�K�K���K K K ����KtK�K�K���K K K ����KaK�K�K���K K K ����KtK�K�K���K K K ����KiK�K�K���K K K ����KwK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KqK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K6K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KtK�K�K���K K K ����KkK�K�K���K K K ����K-K�K�K���K K K ����KaK�K�K���K K K ����KtK�K�K���K K K ����KaK�K�K���K K K ����KsK�K�K���K K K ����KaK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KuK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KBK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KtK�K�K���K K K ����KeK�K�K���K K K ����K-K�K�K���K K K ����KcK�K�K���K K K ����KtK�K�K���K K K ����KcK�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����KdK�K�K���K K K ����K-K�K�K���K K K ����KkK�K�K���K K K ����KaK�K�K���K K K ����KkK�K�K���K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KcK�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KcK�K�K���K K K ����KeK�K�K���K K K ����KfK�K�K���K K K ����KkK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KDK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KgK�K�K���K K K ����KkK�K�K���K K K ����KuK�K�K���K K K ����K-K�K�K���K K K ����KdK�K�K���K K K ����KkK�K�K���K K K ����KdK�K�K���K K K ����KrK�K�K���K K K ����KiK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K7K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KhK�K�K���K K K ����KhK�K�K���K K K ����KeK�K�K���K K K ����KpK�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����KlK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����KdK�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����KZK�K�K���K K K ����KdK�K�K���K K K ����KZK�K�K���K K K ����KiK�K�K���K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KkK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K+K�K�K���K K K ����K-K�K�K���K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����KoK�K�K���K K K ����KdK�K�K���K K K ����KeK�K�K���K K K ����K+K�K�K���K K K ����KLK�K�K���K K K ����K+K�K�K���K K K ����KLK�K�K���K K K ����KLK�K�K���K K K ����KBK�K�K���K K K ����K+K�K�K���K K K ����KSK�K�K���K K K ����KGK�K�K���K K K ����K9K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KKK�K�K���K K K ����K1K�K�K���K K K ����K-K�K�K���K K K ����KmK�K�K���K K K ����KKK�K�K���K K K ����KmK�K�K���K K K ����K!K�K�K���K K K ����KdK�K�K���K K K ����K1K�K�K���K K K ����KoK�K�K���K K K ����K1K�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K1K�K�K���K K K ����KcK�K�K���K K K ����KrK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KCK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����KbK�K�K���K K K ����KyK�K�K���K K K ����KbK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KnK�K�K���K K K ����K K�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KmK�K�K���K K K ����K K�K�K���K K K ����KrK�K�K���K K K ����KeK�K�K���K K K ����KcK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KlK�K�K���K K K ����KIK�K�K���K K K ����K-K�K�K���K K K ����KiK�K�K���K K K ����KlK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����KbK�K�K���K K K ����KLK�K�K���K K K ����KgK�K�K���K K K ����KLK�K�K���K K K ����KgK�K�K���K K K ����KgK�K�K���K K K ����KbK�K�K���K K K ����KIK�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����KeK�K�K���K K K ����KsK�K�K���K K K ����KeK�K�K���K K K ����KsK�K�K���K K K ����KsK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����KnK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KpK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����K K�K�K���K K K ����KoK�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����KwK�K�K���K K K ����KaK�K�K���K K K ����KwK�K�K���K K K ����KwK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KfK�K�K���K K K ����KnK�K�K���K K K ����K-K�K�K���K K K ����KfK�K�K���K K K ����KfK�K�K���K K K ����KfK�K�K���K K K ����K K K K ��K K K ����KKK�K�K���K K K ����KtK�K�K���K K K ����KoK�K�K���K K K ����KtK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K�K�K���K K K ����KHK�K�K���K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����KhK�K�K���K K K ����KrK�K�K���K K K ����KhK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KrK�K�K���K K K ����KHK�K�K���K K K ����K-K�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����KeK�K�K���K K K ����KdK�K�K���K K K ����e(KeK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����KfK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KLK�K�K���K K K ����KBK�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����KbK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K5K�K�K���K K K ����KlK�K�K���K K K ����K-K�K�K���K K K ����K3K�K�K���K K K ����K5K�K�K���K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KlK�K�K���K K K ����KLK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����KmK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KgK�K�K���K K K ����KbK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KhK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KwK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KBK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ���       K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K@KKYK���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K#KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K#KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e��bjP  jP  �width�K#�turn�M��xConst�Kj�}  h�yConst�KF�height�K�MessageHandler��
MessageSys��Messages���)��}�(�messages�]�(�Kyle acquired 19 coins��Kyle picked up Green Herb��'Kyle picked up Scroll of Lightning Bolt��Kyle picked up +1 Iron Helm��Kyle picked up Bomb��Kyle picked up Longsword��Kyle picked up Longsword��Kyle picked up +1 Leather Helm��Zombie dropped Longsword��Zombie dropped +1 Leather Helm��Zombie was killed by Kyle��Zombie is afraid!��Kyle attacked Zombie for 3��Zombie attacked Kyle for 5��Kyle attacked Zombie for 3��Zombie attacked Kyle for 5��Kyle picked up +1 Iron Helm��Zombie attacked Kyle for 5��Skeleton Knight dropped Bomb��!Skeleton Knight dropped Longsword��$Skeleton Knight dropped +1 Iron Helm��"Skeleton Knight was killed by Kyle��Skeleton Knight is afraid!��#Kyle attacked Skeleton Knight for 2��#Skeleton Knight attacked Kyle for 6��Kyle missed Skeleton Knight��#Skeleton Knight attacked Kyle for 6��#Kyle attacked Skeleton Knight for 2��#Skeleton Knight attacked Kyle for 6��#Kyle attacked Skeleton Knight for 2��Skeleton Knight missed Kyle��#Kyle attacked Skeleton Knight for 2��#Skeleton Knight attacked Kyle for 6��Kyle acquired 13 coins��Kyle picked up Longsword��Kyle picked up Chain Shirt��Kyle acquired 6 Arrows��Kyle acquired 9 coins��Kyle picked up Green Herb��Kyle picked up Iron Helm��Kyle picked up Buckler��Kyle picked up Bomb��Kyle acquired 4 coins��Kyle picked up Longsword��Kyle picked up Longsword��Kyle picked up Iron Helm��Skeleton Knight dropped Bomb��!Skeleton Knight dropped Longsword��!Skeleton Knight dropped Iron Helm��"Skeleton Knight was killed by Kyle��Skeleton Knight is afraid!��#Kyle attacked Skeleton Knight for 3��#Skeleton Knight attacked Kyle for 4��#Kyle attacked Skeleton Knight for 3��#Skeleton Knight attacked Kyle for 4��Kyle picked up Iron Helm��#Skeleton Knight attacked Kyle for 4��"Skeleton Knight dropped Gold Coins��!Skeleton Knight dropped Longsword��!Skeleton Knight dropped Iron Helm��"Skeleton Knight was killed by Kyle��Skeleton Knight is afraid!��#Kyle attacked Skeleton Knight for 3��#Skeleton Knight attacked Kyle for 4��#Kyle attacked Skeleton Knight for 3��Kyle waited...��Kyle acquired 7 coins��Kyle picked up Longsword��Kyle picked up Iron Helm��"Skeleton Knight dropped Gold Coins��!Skeleton Knight dropped Longsword��!Skeleton Knight dropped Iron Helm��"Skeleton Knight was killed by Kyle��Skeleton Knight is afraid!��#Kyle attacked Skeleton Knight for 3��#Skeleton Knight attacked Kyle for 4��#Kyle attacked Skeleton Knight for 3��#Skeleton Knight attacked Kyle for 4��Kyle picked up Green Herb��'Kyle picked up Scroll of Lightning Bolt��Kyle picked up Longsword��Kyle picked up Longsword��Kyle picked up Iron Helm��0Skeleton Knight dropped Scroll of Lightning Bolt��!Skeleton Knight dropped Longsword��!Skeleton Knight dropped Iron Helm��"Skeleton Knight was killed by Kyle��Skeleton Knight is afraid!��#Kyle attacked Skeleton Knight for 3��#Skeleton Knight attacked Kyle for 4��#Kyle attacked Skeleton Knight for 3��Kyle acquired 15 coins��Kyle picked up Iron Helm��Kyle picked up Wooden Shield��Kyle picked up Iron Helm��Kyle picked up Leather Helm��Zombie dropped Longsword��Zombie dropped Leather Helm��Zombie was killed by Kyle��Zombie is afraid!��Kyle attacked Zombie for 3��Zombie attacked Kyle for 3��Kyle attacked Zombie for 3��Zombie attacked Kyle for 3��Player Ready: Kyle��
Game Start�e�messageLimit�M��retrieveLimit�Kubub�djikstra_Player_Adj�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKKKKNNNNNNNNNNNKKKKKKKKKKKKKK K!K"K#K$K%NNNNNNNNNNNNNNNNNNNNNNe]�(NNNKKKKKNNNNNNNNNNNKNNNNNNNNNNKK K!K"K#K$K%K&NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKK KNNNNNNNNNNNKNNNNNNNNNNK K!K"K#K$K%K&K'NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKK KK NNNNNNNNNNNKNNNNNNNNNNK!K"K#K$K%K&K'K(NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKK KNNNNNNNNNNNKNNNNNNNNNNNK#K$K%K&K'K(K)NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKKKKKKKK	K
KKKKNNNNNNNNNNNNK%K&K'K(K)K*NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNK'NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNK(NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNK)NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK*NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK+NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK,NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK-NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK	NNNNNNNNNNNNNNNNNNNNNNNNNNK.NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK
KKKNNNNNNNNNNNNNNNNNNNNNNNK/NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK0NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNK+K,K-K.K/K0K1K2K3K4K5K6K7K8NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNK*NNNNNNK3K4K5K6K7K8K9NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNK)NNNNNNK4K5K6K7K8K9K:NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNK(NNNNNNK5K6K7K8K9K:K;NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNK'NNNNNNK6K7K8K9K:K;K<NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKKKKKK K!K"K#K$K%K&NNNNNNK7K8K9K:K;K<K=NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNK8K9K:K;K<K=K>NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNK9K:K;K<K=K>K?NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNK:K;K<K=K>K?K@NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK!NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK"NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK#NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNK'K&K%K$NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKSKTKUKVNNNNNNNNNNNNNNNNNNe]�(NNNNK(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKQKRKSKTKUNNNNNNNNNNNNNNNNNNe]�(NNNNK)NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKOKPKQKRKSKTNNNNNNNNNNNNNNNNNNe]�(NNNNK*K+K,K-K.NNNNNNNNNNNNNNNNNNNNNNNNNNNKNKOKPKQKRKSNNNNNNNNNNNNNNNNNNe]�(NNNNK+K,K-K.K/K0K1K2K3K4K5K6K7K8K9K:NNNNNNNNNNNNNNNNKMKNKOKPKQKRNNNNNNNNNNNNNNNNNNe]�(NNNNK,K-K.K/K0NNNNNNNNNNK;K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQNNNNNNNNNNNNNNNNNNe]�(NNNNK-K.K/K0K1NNNNNNNNNNNNNNNNNNNNNNNNNNNKMKNKOKPKQKRNNNNNNNNNNNNNNNNNNe]�(NNNNK.K/K0K1K2NNNNNNNNNNNNNNNNNNNNNNNNNNNKNKOKPKQKRKSNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKOKPKQKRKSKTNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�djikstra_Player_Away�j�|  h2�1B: Dark Crypt��
messageSys�jש  �SeesMap�]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K ee�inSeed�Jv �textWall��Ornate stone wall
�ubh�ej��  jש  j�}  j�}  �cursor�Kubj�}  hj�}  ]�(hQh�h�h�hrej�}  ]�j�}  ]�(KKej�}  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK6K5K4K3K2NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK5K4K3K2K1NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK4K3K2K1K0NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK3K2K1K0K/NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK2K1K0K/K.NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KNNNNNNNNNNNNK
K	KKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK2K1K0K/K.NNNNNNNNNNNNNKNNNNNNNNNNNNK	KKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK3K2K1K0K/NNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK2K1K0NNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK3K2K1NNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKKK KKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK4NNNNNNNNNNNNNNNKNNNNNNNNNNNNNKNNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK5NNNNNNNNNNNNNNNKNNNNNNNNNNNNKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK6NNNNNNNNNNNNNNNKNNNNNNNNNNNNK	KKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK7NNNNNNNNNNNNNNNKKKKKKKKKKKKKK
K	KKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK8NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK	NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK<K;K:K9NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK
NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK=NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK?NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK@NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKANNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKBNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKGKFKEKDKCNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKFKEKDKCKBNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKEKDKCKBKANNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKDKCKBKAK@NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKCKBKAK@K?NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKBKAK@K?K>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKAK@K?K>K=NNNNNNNNNNNNNNNK)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNK>K=K<NNNNNNNNNNNNNNNK*NNNNNNNNNNNNNNNNNKKKKKKK NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNK=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+NNNNNNNNNNNNNNNNNNKKKKK K!NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej�}  j�}  jG�  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNN��I      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK5K4K3K2K1NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK4K3K2K1K0NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK3K2K1K0K/NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK2K1K0K/K.NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK1K0K/K.K-NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKNNNNNNNNNNNNK	KKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK1K0K/K.K-NNNNNNNNNNNNNKNNNNNNNNNNNNKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK2K1K0K/K.NNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK1K0K/NNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKKK KKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK2K1K0NNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKK KK KKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK3NNNNNNNNNNNNNNNKNNNNNNNNNNNNNKNNKKK KKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK4NNNNNNNNNNNNNNNKNNNNNNNNNNNNKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK5NNNNNNNNNNNNNNNKNNNNNNNNNNNNKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK6NNNNNNNNNNNNNNNKKKKKKKKKKKKK
K	KKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK7NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK;K:K9K8NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK	NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK<NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK
NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK=NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK?NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK@NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKANNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKBNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKFKEKDKCKBNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKEKDKCKBKANNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKDKCKBKAK@NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKCKBKAK@K?NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKBKAK@K?K>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKAK@K?K>K=NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK@K?K>K=K<NNNNNNNNNNNNNNNK(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNK=K<K;NNNNNNNNNNNNNNNK)NNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNK<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*NNNNNNNNNNNNNNNNNNKKKKKK NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej��  j
O  h2�2B: Dark Crypt�j��  jש  j��  ]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K KK K KKKKKKKKK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K KK K KKKKKKKKK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K eejƪ  M�jǪ  jȪ  ubh/h�j  K7j  KEj  Kh�hh2h ub�skillPoints�Kj0  ]�hHKj/  Kdh-]�(KKYK�eh2�Kyle�ub.