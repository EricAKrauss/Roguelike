��      �__main__��Game���)��}�(�loadRequest���console��tdl��Console���)��KYK*]�(K K K K ��K K K ����KKK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KLK�K�K���K K K ����KEK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KRK�K�K���K K K ����KPK�K�K���K K K ����KAK�K�K���K K K ����K K K K ��K K K ����KAK�K�K���K K K ����KWK�K�K���K K K ����K K K K ��K K K ����KGK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KSK�K�K���K K K ����KSK�K�K���K K K ����KZK�K�K���K K K ����KKK�K�K���K K K ����K-K�K�K���K K K ����KKK�K�K���K K K ����KZK�K�K���K K K ����KKK�K�K���K K K ����KZK�K�K���K K K ����KZK�K�K���K K K ����KZK�K�K���K K K ����KZK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KxK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KaK�K�K���K K K ����KoK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KoK�K�K���K K K ����KyK�K�K���K K K ����K-K�K�K���K K K ����KyK�K�K���K K K ����KoK�K�K���K K K ����KyK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����KyK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����KFK�K�K���K K K ����K K K K ��K K K ����KvK�K�K���K K K ����KpK�K�K���K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KnK�K�K���K K K ����KwK�K�K���K K K ����KmK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KmK�K�K���K K K ����KlK�K�K���K K K ����K-K�K�K���K K K ����KlK�K�K���K K K ����KmK�K�K���K K K ����KlK�K�K���K K K ����KmK�K�K���K K K ����KmK�K�K���K K K ����KmK�K�K���K K K ����KmK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KgK�K�K���K K K ����K K K K ��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KlK�K�K���K K K ����KlK�K�K���K K K ����KbK�K�K���K K K ����KeK�K�K���K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KbK�K�K���K K K ����KeK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KbK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����KwK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KhK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KiK�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����KiK�K�K���K K K ����K K�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K3K�K�K���K K K ����K K K K ��K K K ����KhK�K�K���K K K ����K K K K ��K K K ����KsK�K�K���K K K ����K:K�K�K���K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����KeK�K�K���K K K ����KpK�K�K���K K K ����K-K�K�K���K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����KaK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KPK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K6K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����KiK�K�K���K K K ����K-K�K�K���K K K ����KtK�K�K���K K K ����K K�K�K���K K K ����KtK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KcK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K1K�K�K���K K K ����K4K�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K7K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����KcK�K�K���K K K ����K-K�K�K���K K K ����KtK�K�K���K K K ����KaK�K�K���K K K ����KtK�K�K���K K K ����KiK�K�K���K K K ����KwK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KcK�K�K���K K K ����KqK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K6K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KtK�K�K���K K K ����KkK�K�K���K K K ����K-K�K�K���K K K ����KaK�K�K���K K K ����KtK�K�K���K K K ����KaK�K�K���K K K ����KsK�K�K���K K K ����KaK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KkK�K�K���K K K ����KuK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KBK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KKK�K�K���K K K ����KKK�K�K���K K K ����KtK�K�K���K K K ����KeK�K�K���K K K ����K-K�K�K���K K K ����KcK�K�K���K K K ����KtK�K�K���K K K ����KcK�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K:K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K0K�K�K���K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KaK�K�K���K K K ����KdK�K�K���K K K ����K-K�K�K���K K K ����KkK�K�K���K K K ����KaK�K�K���K K K ����KkK�K�K���K K K ����KaK�K�K���K K K ����K K�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K/K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����KiK�K�K���K K K ����KcK�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KcK�K�K���K K K ����KeK�K�K���K K K ����KfK�K�K���K K K ����KkK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KDK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K2K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����KgK�K�K���K K K ����KkK�K�K���K K K ����KuK�K�K���K K K ����K-K�K�K���K K K ����KdK�K�K���K K K ����KkK�K�K���K K K ����KdK�K�K���K K K ����KrK�K�K���K K K ����KiK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KuK�K�K���K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KaK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K7K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KhK�K�K���K K K ����KhK�K�K���K K K ����KeK�K�K���K K K ����KpK�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����KlK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K5K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����KtK�K�K���K K K ����KdK�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����KZK�K�K���K K K ����KdK�K�K���K K K ����KZK�K�K���K K K ����KiK�K�K���K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K1K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KkK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K+K�K�K���K K K ����K-K�K�K���K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����KoK�K�K���K K K ����KdK�K�K���K K K ����KeK�K�K���K K K ����K+K�K�K���K K K ����KLK�K�K���K K K ����K+K�K�K���K K K ����KLK�K�K���K K K ����KLK�K�K���K K K ����KBK�K�K���K K K ����K+K�K�K���K K K ����KSK�K�K���K K K ����KGK�K�K���K K K ����K9K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KKK�K�K���K K K ����K1K�K�K���K K K ����K-K�K�K���K K K ����KmK�K�K���K K K ����KKK�K�K���K K K ����KmK�K�K���K K K ����K!K�K�K���K K K ����KdK�K�K���K K K ����K1K�K�K���K K K ����KoK�K�K���K K K ����K1K�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K1K�K�K���K K K ����KcK�K�K���K K K ����KrK�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KCK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KyK�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����KbK�K�K���K K K ����KyK�K�K���K K K ����KbK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KnK�K�K���K K K ����K K�K�K���K K K ����KnK�K�K���K K K ����KnK�K�K���K K K ����KmK�K�K���K K K ����K K�K�K���K K K ����KrK�K�K���K K K ����KeK�K�K���K K K ����KcK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KlK�K�K���K K K ����KIK�K�K���K K K ����K-K�K�K���K K K ����KiK�K�K���K K K ����KlK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����KbK�K�K���K K K ����KLK�K�K���K K K ����KgK�K�K���K K K ����KLK�K�K���K K K ����KgK�K�K���K K K ����KgK�K�K���K K K ����KbK�K�K���K K K ����KIK�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KyK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����K-K�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����KeK�K�K���K K K ����KsK�K�K���K K K ����KeK�K�K���K K K ����KsK�K�K���K K K ����KsK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����KlK�K�K���K K K ����KnK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KpK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KpK�K�K���K K K ����KpK�K�K���K K K ����K K�K�K���K K K ����KoK�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KaK�K�K���K K K ����KwK�K�K���K K K ����KaK�K�K���K K K ����KwK�K�K���K K K ����KwK�K�K���K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KlK�K�K���K K K ����K K�K�K���K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KeK�K�K���K K K ����KfK�K�K���K K K ����KnK�K�K���K K K ����K-K�K�K���K K K ����KfK�K�K���K K K ����KfK�K�K���K K K ����KfK�K�K���K K K ����K K K K ��K K K ����KKK�K�K���K K K ����KtK�K�K���K K K ����KoK�K�K���K K K ����KtK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K�K�K���K K K ����KHK�K�K���K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����KoK�K�K���K K K ����K K�K�K���K K K ����K-K�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����KyK�K�K���K K K ����KhK�K�K���K K K ����KrK�K�K���K K K ����KhK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����KoK�K�K���K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KrK�K�K���K K K ����KHK�K�K���K K K ����K-K�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����KeK�K�K���K K K ����KdK�K�K���K K K ����e(KeK�K�K���K K K ����KdK�K�K���K K K ����KdK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����KfK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KLK�K�K���K K K ����KBK�K�K���K K K ����K K�K�K���K K K ����KeK�K�K���K K K ����K-K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����KrK�K�K���K K K ����K K K K ��K K K ����KrK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K�K�K���K K K ����KbK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����KoK�K�K���K K K ����K5K�K�K���K K K ����KlK�K�K���K K K ����K-K�K�K���K K K ����K3K�K�K���K K K ����K5K�K�K���K K K ����K3K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KlK�K�K���K K K ����KLK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����KmK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KHK�K�K���K K K ����K K K K ��K K K ����KHK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KgK�K�K���K K K ����KbK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����KeK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KsK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KhK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KwK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KmK�K�K���K K K ����K K K K ��K K K ����KmK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����K K�K�K���K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KiK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����KdK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KnK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KgK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KBK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KoK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KlK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K.K�K�K���K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����KtK�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K@KKYK���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K#KdKdKd��K K K ����K#K|K�K��K K K ����K.K�K�K���K K K ����K#K|K�K��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K.KdKdKd��K K K ����K.K�K�K���K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K#KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K#KdKdKd��K K K ����K.KdKdKd��K K K ����K#KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K KdKdKd��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K|K�K�K���K K K ����K-K�K�K���K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e(K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K �      K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����K K K K ��K K K ����e��b�	levelList��LevelManager�j�+  ��)��}�(�nextSeed�M&j�+  ]�(�LevelTypes.LevelTypes��Crypt���)��}�(�cLevel�K�args�]�(KKKKKKe�itemList�]�(�Items.Consumables��	GreenHerb���j�+  �Bundle_Of_Arrows���j�+  �	Time_Bomb���j�+  �Scroll_of_Fireball���j�+  �Scroll_of_Lightning_Bolt����Items.Weapons��Staff���j�+  �Iron_Shield���j�+  �Buckler���j�+  �Wooden_Shield���j�+  �	Longsword���j�+  �
Greatsword���j�+  �Bow���j�+  �Spear���j�+  �Dagger����Items.Armors��Cloth_Shirt���j
,  �	Cloth_Hat���j
,  �Leather_Shirt���j
,  �Leather_Helm���j
,  �Iron_Breastplate���j
,  �	Iron_Helm���j
,  �Chain_Shirt���j
,  �
Chain_Helm���e�healingList�]�j�+  a�	equipList�]�(j�+  j�+  j�+  j�+  j,  j,  j,  j,  j	,  j,  j,  j,  j,  j,  j,  j,  j,  e�stairsUp�]�(KKe�	eliteList�]��Enemies.Undead��Cultist���a�Objects�}�(K �Object�j(,  ��)��}�(�pLevel�j�+  �char��*��ID�K �row�K�col�Kj(,  �LevelTypes.Decorations��Ritual_Circle���)��}�(�name��Ritual Circle��pObject�j*,  j-,  j.,  ubj7,  j8,  ubKj),  )��}�(j,,  j�+  j-,  �~�j/,  Kj0,  Kj1,  Kj(,  �Features.Features��Brush���)��}�(j9,  j:,  �color�]�(KKnKej-,  j<,  j7,  j>,  ubj7,  j>,  ubKj),  )��}�(j,,  j�+  j-,  �+�j/,  Kj0,  Kj1,  K"j(,  j�+  )��}�(�
equippable���
consumable���healNum�Kj9,  jD,  �type�jJ,  jB,  ]�(K�K�K�ej-,  jF,  j7,  �
Green Herb�ubj7,  �Health�ubKj),  )��}�(j,,  j�+  j-,  j<,  j/,  Kj0,  Kj1,  Kj(,  j?,  )��}�(j9,  jP,  jB,  jC,  j-,  j<,  j7,  j>,  ubj7,  j>,  ubKj),  )��}�(j,,  j�+  j-,  �=�j/,  Kj0,  Kj1,  Kj(,  j=,  �Chest���)��}�(�items�]�(j�+  )��}�(�
arrowCount�KjJ,  �jL,  jJ,  jB,  jM,  j-,  �i�jI,  �j7,  �Bundle of Arrows�ubj�+  )��}�(�level�KjI,  �jJ,  ��spell��	Abilities��Fireball���jL,  �scroll�jB,  jM,  j-,  �s�j7,  �Scroll of Fireball�ubj,  )��}�(�armorVal�Kjd,  KjI,  �jJ,  ��weight�KjL,  �armor�jB,  jM,  j-,  �?��	throwable��j7,  �Leather Shirt�ubj�+  �
Gold_Coins���)��}�(jI,  �jJ,  �jL,  jJ,  jB,  ]�(K�K�Kej-,  �$��coins�K	j7,  �
Gold Coins�ubej9,  jT,  jB,  ]�(KQKOKej-,  jV,  j7,  jW,  ubj7,  jW,  ubKj),  )��}�(j,,  j�+  j-,  �x�j/,  Kj0,  Kj1,  K j(,  j#,  �Skeleton_Knight���)��}�(jd,  K�exp�K j-,  j,  �
dropChance�K(�
alliesList�]�(j},  j),  )��}�(j,,  j�+  j-,  j,  j/,  K	j0,  Kj1,  K%j(,  j#,  �Zombie���)��}�(jd,  Kj�,  K j-,  j,  j�,  K(j�,  ]�(j},  j�,  e�power�K�playerControlled���helmet�j,  )��}�(jn,  K
jd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �Leather Helm�ub�armorPen�K �gold�K�
healthTemp�K �dodge�K �	sightDist�K	�
initiative�K�health�K�leftHand�N�	cowardice�G        �canMove���
countering��j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  js,  ub�range�K�visible���	rightRing�N�accuracy�K �necklace�N�	rightHand�j,  )��}�(jd,  Kj-,  jq,  jL,  �1H�jI,  �jJ,  ��addPower��j�,  Kj�,  Kjo,  K�magPower�K�
usesArrows��jB,  jM,  j�,  Kjr,  �j7,  j ,  ub�lastPlayerLoc�Njn,  K �isAfraid���blocking���arrows�K �lastPlayerMap�N�	healthMax�K�hearingDist�K�leftRing�N�invertColor���
hitEffects�]�j9,  j�,  �expNext�Kd�effects�]��
stealthVal�K jB,  ]�(K�KKej7,  j�,  ubj7,  �Enemy�ubej�,  Kj�,  �j�,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �	Iron Helm�ubj�,  K j�,  Kj�,  K j�,  K j�,  Kj�,  Kj�,  Kj�,  j�+  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �jn,  Kj�,  K jo,  Kj�,  K jB,  jM,  j�,  Kj�,  �jr,  �j7,  �Wooden Shield�ubj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  js,  ubj�,  Kj�,  �j�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  Kjr,  �j7,  j ,  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  j},  j�,  Kdj�,  ]�j�,  K jB,  j�,  j7,  �Skeleton Knight�ubj7,  j�,  ubKj),  )��}�(j,,  j�+  j-,  �S�j/,  Kj0,  Kj1,  Kj(,  �Features.Stairs��StairUp���)��}�(j9,  j�,  j,,  j�+  �moveCost�Kj/,  J����j0,  Kj1,  Kj(,  Nj7,  �Stairs�ubj7,  �	Stairs Up�ubKj),  )��}�(j,,  j�+  j-,  �@�j/,  Kj0,  K(j1,  K)j(,  �Player�j�,  ��)��}�(jd,  Kj�,  K#�recalcTimer�K �skills�}�(�3�jh,  �4�jf,  �Lightning_Bolt����7�jf,  �Ready_for_Battle����5�jf,  �Block����6�jf,  �Rending_Blow����1�jf,  �Charge����2�jf,  �Shocking_Grasp���u�
prevTarget�Nj�,  Kj�,  �j�,  j,  )��}�(jn,  K
jd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  j�,  ubj�,  K j�,  KCj�,  K j�,  K j�,  Kj�,  Kjp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �Cloth Shirt�ubj�,  j�+  �Tome���)��}�(jd,  Kj-,  jq,  jL,  �0H�jI,  �jJ,  �j�,  �j�,  Kj�,  K jo,  Kj�,  Kj�,  �jB,  jM,  j�,  K jr,  �j7,  j�,  ubj�,  �j�,  �j[,  ]�(j�+  )��}�(jI,  �jJ,  �jK,  KjL,  jJ,  jB,  jM,  j-,  jF,  j7,  jN,  ubj�+  )��}�(jI,  �jJ,  �jK,  KjL,  jJ,  jB,  jM,  j-,  jF,  j7,  jN,  ubj,  )��}�(jn,  K
jd,  KjI,  �jJ,  �jo,  Kj9,  NjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  j�,  ubj,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  j�,  ubj�+  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �jn,  Kj�,  K jo,  Kj�,  K jB,  jM,  j�,  Kj�,  �jr,  �j7,  j�,  ubj,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  j�,  ubj,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  Kj9,  NjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  j�,  ubj,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j9,  Nj�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  Kjr,  �j7,  j ,  ubj,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j9,  Nj�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  Kjr,  �j7,  j ,  ubj�+  )��}�(jd,  KjI,  �jJ,  �je,  j�,  j9,  NjL,  ji,  jB,  jM,  j-,  jj,  j7,  �Scroll of Lightning Bolt�ubj�+  )��}�(jI,  �jJ,  �jK,  Kj9,  NjL,  jJ,  jB,  jM,  j-,  jF,  j7,  jN,  ubj,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  Kj9,  NjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  j�,  ubj,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j9,  Nj�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  Kjr,  �j7,  j ,  ubj,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  Kj9,  NjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  j�,  ubj,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  Kj9,  NjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  j�,  ubj,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j9,  Nj�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  Kjr,  �j7,  j ,  ubj,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j9,  Nj�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  Kjr,  �j7,  j ,  ubj�+  )��}�(jd,  Kj-,  �o�jL,  jJ,  jI,  �jJ,  �j9,  N�dur�KjB,  jM,  j�,  K j7,  �Bomb��desc��Explodes up after 3 turns��damage�K�radius�Kubj�+  )��}�(jd,  Kj-,  jq,  jL,  j -  jI,  �jJ,  �j�,  �jn,  Kj�,  K jo,  Kj�,  K jB,  jM,  j�,  Kj�,  �jr,  �j7,  j�+  ubj,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  j�,  ubj�+  )��}�(jI,  �jJ,  �jK,  KjL,  jJ,  jB,  jM,  j-,  jF,  j7,  jN,  ubj,  )��}�(jn,  K#jd,  KjI,  �jJ,  �jo,  K#jL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �Chain Shirt�ubj,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  Kjr,  �j7,  j ,  ubj,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  Kj9,  NjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Iron Helm�ubj,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  Kj9,  NjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Helm�ubj,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j9,  Nj�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j ,  ubj,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j9,  Nj�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j ,  ubj�+  )��}�(jd,  Kj-,  j'-  jL,  jJ,  jI,  �jJ,  �j9,  Nj(-  KjB,  jM,  j�,  K j7,  j)-  j*-  j+-  j,-  Kj--  Kubj,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Iron Helm�ubj�+  )��}�(jd,  KjI,  �jJ,  �je,  j�,  jL,  ji,  jB,  jM,  j-,  jj,  j7,  j-  ubj�+  )��}�(jI,  �jJ,  �jK,  K jL,  jJ,  jB,  jM,  j-,  jF,  j7,  jN,  ubej�,  K�j�,  ��
baseHealth�Mj�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  �2H�jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  Kjr,  �j7,  j,  ubj-,  j�,  jn,  K �
leftScroll�Nj�,  �j�,  K�Class��Player_Classes��
Spellsword���j�,  Mj�,  N�	recalcMax�K �healthCurve�G?�333333�rightScroll�Nj�,  �j�,  ]��skillLevels�}�(j�,  K j�,  K j�,  K j�,  K j�,  K j�,  K j�,  K uj9,  j),  )��}�(j,,  j�+  )��}�(j�+  Kj�+  ]�(KKKKKKej�+  ]�(j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  j�+  j,  j,  j,  j,  j	,  j,  j,  j,  j,  j,  j,  j,  j,  ej,  ]�j�+  aj,  ]�(j�+  j�+  j�+  j�+  j,  j,  j,  j,  j	,  j,  j,  j,  j,  j,  j,  j,  j,  ej,  ]�(K/K/ej!,  j",  j&,  }�(K@j),  )��}�(j,,  j]-  j-,  jq,  j/,  K@j0,  K>j1,  K
j(,  j�+  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j9,  je-  jn,  Kj�,  K jo,  Kj�,  K jB,  jM,  j�,  Kj�,  �jr,  �j7,  j�,  ubj7,  �Item�ubKCj),  )��}�(j,,  j]-  j-,  j,  j/,  KCj0,  K?j1,  K	j(,  j�,  )��}�(jd,  Kj�,  K j-,  j,  j�,  K(j�,  ]�(jj-  j),  )��}�(j,,  j]-  j-,  j,  j/,  KDj0,  K@j1,  K
j(,  j�,  )��}�(jd,  Kj�,  K j-,  j,  j�,  K(j�,  ]�(jj-  jo-  j),  )��}�(j,,  j]-  j-,  j,  j/,  KFj0,  KBj1,  K
j(,  j�,  )��}�(jd,  Kj�,  K j-,  j,  j�,  K(j�,  ]�(jj-  jo-  jt-  ej�,  Kj�,  �j�,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Helm�ubj�,  K j�,  Kj�,  K j�,  K j�,  K	j�,  Kj�,  Kj�,  Nj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Shirt�ubj�,  Kj�,  �j�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j ,  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  jt-  j�,  Kdj�,  ]�j�,  K jB,  j�,  j7,  j�,  ubj7,  j�,  ubej�,  Kj�,  �j�,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Helm�ubj�,  K j�,  K
j�,  K j�,  K j�,  K	j�,  Kj�,  Kj�,  Nj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Shirt�ubj�,  Kj�,  �j�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j ,  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  jo-  j�,  Kdj�,  ]�j�,  K jB,  j�,  j7,  j�,  ubj7,  j�,  ubjt-  ej�,  Kj�,  �j�,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Helm�ubj�,  K j�,  Kj�,  K j�,  K j�,  K	j�,  Kj�,  Kj�,  Nj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Shirt�ubj�,  Kj�,  �j�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j ,  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  jj-  j�,  Kdj�,  ]�j�,  K jB,  j�,  j7,  j�,  ubj7,  j�,  ubKDjo-  KEj),  )��}�(j,,  j]-  j-,  jV,  j/,  KEj0,  KAj1,  K2j(,  jX,  )��}�(j[,  ]�j9,  j�-  jB,  jM,  j-,  jV,  j7,  jW,  ubj7,  jW,  ubKFjt-  KGj),  )��}�(j,,  j]-  j-,  jV,  j/,  KGj0,  KCj1,  K
j(,  jX,  )��}�(j[,  ]�(j,  )��}�(jd,  Kj-,  jq,  jL,  jO-  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j,  ubj,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  K
jL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Chain Helm�ubj,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Cloth Hat�ubju,  )��}�(jI,  �jJ,  �jL,  jJ,  jB,  jx,  j-,  jy,  jz,  Kj7,  j{,  ubej9,  j�-  jB,  j|,  j-,  jV,  j7,  jW,  ubj7,  jW,  ubKHj),  )��}�(j,,  j]-  j-,  j.,  j/,  KHj0,  KDj1,  K,j(,  j2,  �Altar���)��}�(j7,  j�-  j9,  j�-  j-,  j.,  ubj7,  j�-  ubKIj),  )��}�(j,,  j]-  j-,  jq,  j/,  KIj0,  K<j1,  K+j(,  j9-  j7,  j;-  ubKJj),  )��}�(j,,  j]-  j-,  jq,  j/,  KJj0,  K<j1,  K+j(,  j?-  j7,  j ,  ubKKj),  )��}�(j,,  j]-  j-,  j'-  j/,  KKj0,  K<j1,  K+j(,  jC-  j7,  j)-  ubKLj),  )��}�(j,,  j]-  j-,  jq,  j/,  KLj0,  K<j1,  K,j(,  j<-  j7,  j>-  ubKMj),  )��}�(j,,  j]-  j-,  jq,  j/,  KMj0,  K<j1,  K,j(,  jA-  j7,  j ,  ubK%j),  )��}�(j,,  j]-  j-,  �E�j/,  K%j0,  Kj1,  Kj(,  j�,  �	StairDown���)��}�(j,,  j]-  j9,  j�-  j/,  J����j0,  Kj�,  Kj(,  Nj1,  Kj7,  j�,  ubj7,  �Stairs Down�ubK&j),  )��}�(j,,  j]-  j-,  j.,  j/,  K&j0,  Kj1,  Kj(,  j4,  )��}�(j7,  j8,  j9,  j�-  j-,  j.,  ubj7,  j8,  ubK'j),  )��}�(j,,  j]-  j-,  j,  j/,  K'j0,  Kj1,  Kj(,  j�,  )��}�(jd,  Kj�,  K j-,  j,  j�,  K(j�,  ]�(j�-  j),  )��}�(j,,  j]-  j-,  j,  j/,  K(j0,  Kj1,  Kj(,  j�,  )��}�(jd,  Kj�,  K j-,  j,  j�,  K(j�,  ]�(j�-  j�-  j),  )��}�(j,,  j]-  j-,  �X�j/,  K)j0,  Kj1,  Kj(,  j%,  )��}�(jd,  Kj�,  K j-,  j�-  j�,  K(j�,  ]�(j�-  j�-  j�-  ej�,  Kj�,  �j�,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Cloth Hat�ubj�,  K j�,  Kj�,  K j�,  K j�,  Kj�,  Kj�,  Kj�,  j�,  )��}�(jd,  Kj-,  jq,  jL,  j -  jI,  �jJ,  �j�,  �j�,  Kj�,  K jo,  Kj�,  Kj�,  �jB,  jM,  j�,  K jr,  �j7,  j�,  ubj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Cloth Shirt�ubj�,  Kj�,  �j�,  Nj�,  K �cdMax�Kj�,  Nj�,  j�+  )��}�(jd,  Kj-,  jq,  jL,  jO-  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j�+  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  j�-  j�,  Kdj�,  ]�j�,  K jK,  K jB,  j�,  �cd�Kpj7,  �Robed Cultist�ubj7,  j�,  ubej�,  Kj�,  �j�,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Iron Helm�ubj�,  K j�,  Kj�,  K j�,  K j�,  Kj�,  Kj�,  Kj�,  j�+  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �jn,  Kj�,  K jo,  Kj�,  K jB,  jM,  j�,  Kj�,  �jr,  �j7,  j�,  ubj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Shirt�ubj�,  Kj�,  �j�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j ,  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  j�-  j�,  Kdj�,  ]�j�,  K jB,  j�,  j7,  j�,  ubj7,  j�,  ubj�-  ej�,  Kj�,  �j�,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Iron Helm�ubj�,  K j�,  Kj�,  K j�,  K j�,  Kj�,  Kj�,  Kj�,  j�+  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �jn,  Kj�,  K jo,  Kj�,  K jB,  jM,  j�,  Kj�,  �jr,  �j7,  j�,  ubj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Shirt�ubj�,  Kj�,  �j�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j ,  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  j�-  j�,  Kdj�,  ]�j�,  K jB,  j�,  j7,  j�,  ubj7,  j�,  ubK(j�-  K)j�-  K*j),  )��}�(j,,  j]-  j-,  j,  j/,  K*j0,  Kj1,  K-j(,  j�,  )��}�(jd,  Kj�,  K j-,  j,  j�,  K(j�,  ]�j.  aj�,  Kj�,  �j�,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Helm�ubj�,  K j�,  K	j�,  K j�,  K j�,  K	j�,  Kj�,  Kj�,  Nj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Shirt�ubj�,  Kj�,  �j�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j ,  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  j.  j�,  Kdj�,  ]�j�,  K jB,  j�,  j7,  j�,  ubj7,  j�,  ubK+j),  )��}�(j,,  j]-  j-,  j,  j/,  K+j0,  Kj1,  Kj(,  j�,  )��}�(jd,  Kj�,  K j-,  j,  j�,  K(j�,  ]�(j.  j),  )��}�(j,,  j]-  j-,  j,  j/,  K4j0,  Kj1,  Kj(,  j�,  )��}�(jd,  Kj�,  K j-,  j,  j�,  K(j�,  ]�(j.  j.  ej�,  Kj�,  �j�,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Iron Helm�ubj�,  K j�,  Kj�,  K j�,  K j�,  Kj�,  Kj�,  Kj�,  j�+  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �jn,  Kj�,  K jo,  Kj�,  K jB,  jM,  j�,  Kj�,  �jr,  �j7,  j�,  ubj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Shirt�ubj�,  Kj�,  �j�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j ,  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  j.  j�,  Kdj�,  ]�j�,  K jB,  j�,  j7,  j�,  ubj7,  j�,  ubej�,  Kj�,  �j�,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Helm�ubj�,  K j�,  Kj�,  K j�,  K j�,  K	j�,  Kj�,  Kj�,  Nj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Shirt�ubj�,  Kj�,  �j�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j ,  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  j.  j�,  Kdj�,  ]�j�,  K jB,  j�,  j7,  j�,  ubj7,  j�,  ubK,j),  )��}�(j,,  j]-  j-,  j.,  j/,  K,j0,  Kj1,  K,j(,  j�-  )��}�(j7,  j�-  j9,  j6.  j-,  j.,  ubj7,  j�-  ubK-j),  )��}�(j,,  j]-  j-,  j.,  j/,  K-j0,  Kj1,  K-j(,  j4,  )��}�(j7,  j8,  j9,  j:.  j-,  j.,  ubj7,  j8,  ubK.j),  )��}�(j,,  j]-  j-,  j.,  j/,  K.j0,  Kj1,  K,j(,  j2,  �Pile_of_Bones���)��}�(j7,  �Pile of Bones�j9,  j>.  j-,  j.,  ubj7,  jD.  ubK/j),  )��}�(j,,  j]-  j-,  j.,  j/,  K/j0,  Kj1,  K-j(,  j�-  )��}�(j7,  j�-  j9,  jE.  j-,  j.,  ubj7,  j�-  ubK0j),  )��}�(j,,  j]-  j-,  jF,  j/,  K0j0,  Kj1,  K
j(,  j�+  )��}�(jI,  �jJ,  �jK,  K j9,  jI.  jL,  jJ,  jB,  jM,  j-,  jF,  j7,  jN,  ubj7,  jO,  ubK1j),  )��}�(j,,  j]-  j-,  j.,  j/,  K1j0,  Kj1,  K,j(,  j�-  )��}�(j7,  j�-  j9,  jM.  j-,  j.,  ubj7,  j�-  ubK2j),  )��}�(j,,  j]-  j-,  j.,  j/,  K2j0,  Kj1,  K-j(,  j4,  )��}�(j7,  j8,  j9,  jQ.  j-,  j.,  ubj7,  j8,  ubK3j),  )��}�(j,,  j]-  j-,  j�-  j/,  K3j0,  Kj1,  K1j(,  j%,  )��}�(jd,  Kj�,  K j-,  j�-  j�,  K(j�,  ]�jU.  aj�,  Kj�,  �j�,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Cloth Hat�ubj�,  K j�,  Kj�,  K j�,  K j�,  Kj�,  Kj�,  Kj�,  j�,  )��}�(jd,  Kj-,  jq,  jL,  j -  jI,  �jJ,  �j�,  �j�,  Kj�,  K jo,  Kj�,  Kj�,  �jB,  jM,  j�,  K jr,  �j7,  j�,  ubj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Cloth Shirt�ubj�,  Kj�,  �j�,  Nj�,  K j�-  Kj�,  Nj�,  j�+  )��}�(jd,  Kj-,  jq,  jL,  jO-  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j�+  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  jU.  j�,  Kdj�,  ]�j�,  K jK,  K jB,  j�,  j�-  Kpj7,  j�-  ubj7,  j�,  ubK4j.  K5j),  )��}�(j,,  j]-  j-,  j,  j/,  K5j0,  K&j1,  Kj(,  j�,  )��}�(jd,  Kj�,  K j-,  j,  j�,  K(j�,  ]�jg.  aj�,  Kj�,  �j�,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Helm�ubj�,  K j�,  Kj�,  K j�,  K j�,  K	j�,  Kj�,  Kj�,  Nj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  �+1 Leather Shirt�ubj�,  Kj�,  �j�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  K
jr,  �j7,  j ,  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  jg.  j�,  Kdj�,  ]�j�,  K jB,  j�,  j7,  j�,  ubj7,  j�,  ubK6j),  )��}�(j,,  j]-  j-,  j�,  j/,  K6j0,  K/j1,  K/j(,  j�,  )��}�(j9,  jw.  j,,  j]-  j�,  Kj/,  J����j0,  K/j1,  K/j(,  Nj7,  j�,  ubj7,  j�,  ubK7j[-  K8j),  )��}�(j,,  j]-  j-,  j.,  j/,  K8j0,  K0j1,  K*j(,  j4,  )��}�(j7,  j8,  j9,  j{.  j-,  j.,  ubj7,  j8,  ubK9j),  )��}�(j,,  j]-  j-,  j<,  j/,  K9j0,  K4j1,  Kj(,  j?,  )��}�(j9,  j.  jB,  jC,  j-,  j<,  j7,  j>,  ubj7,  j>,  ubK:j),  )��}�(j,,  j]-  j-,  j<,  j/,  K:j0,  K5j1,  K	j(,  j?,  )��}�(j9,  j�.  jB,  jC,  j-,  j<,  j7,  j>,  ubj7,  j>,  ubK;j),  )��}�(j,,  j]-  j-,  j<,  j/,  K;j0,  K5j1,  K
j(,  j?,  )��}�(j9,  j�.  jB,  jC,  j-,  j<,  j7,  j>,  ubj7,  j>,  ubK<j),  )��}�(j,,  j]-  j-,  j<,  j/,  K<j0,  K5j1,  Kj(,  j?,  )��}�(j9,  j�.  jB,  jC,  j-,  j<,  j7,  j>,  ubj7,  j>,  ubK=j),  )��}�(j,,  j]-  j-,  j<,  j/,  K=j0,  K5j1,  Kj(,  j?,  )��}�(j9,  j�.  jB,  jC,  j-,  j<,  j7,  j>,  ubj7,  j>,  ubK>j),  )��}�(j,,  j]-  j-,  j<,  j/,  K>j0,  K6j1,  K	j(,  j?,  )��}�(j9,  j�.  jB,  jC,  j-,  j<,  j7,  j>,  ubj7,  j>,  ubK?j),  )��}�(j,,  j]-  j-,  jF,  j/,  K?j0,  K=j1,  K	j(,  j�+  )��}�(jI,  �jJ,  �jK,  K j9,  j�.  jL,  jJ,  jB,  jM,  j-,  jF,  j7,  jN,  ubj7,  jO,  ubu�CollisionMap�]�(]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKK K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKK KKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKK K K K K KKKKKKKKKKKKKK KKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK K K KKKKKKKKKKKKKK KKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK K K KKKKKKKKKKKKKK KKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK KKKKKKKKKKKKKKKK KKKKKKKKKKKKKK KKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK KKKKKKKKKKKKKKKK KKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK KKKKKKKKKKKKKKKK KKKKKKKKKKKKK K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK KKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K K KKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKK K K KKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKK K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKee�djikstra_Stairs_Down�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKKK KKKKKKKKK	K
KKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNKKKKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNK0K1K2K3K4K5K6NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNK/K0K1K2K3K4K5NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK	KKKKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNK.K/K0K1K2K3K4NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK
K	KKKNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNK-K.K/K0K1K2K3NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNKKKKKKKKKK K!K"K#K$K%K&K'K(K)K*K+K,K-K.K/K0K1K2NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK-K.K/K0K1K2K3NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK.K/K0K1K2K3K4NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK5NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK6NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK7NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK:K9K8NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK;NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK<NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK=NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKkKjKiKhKgKfKeNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKjKiKhKgKfKeKdKcKbKaK`K_K^K]K\K[KZKYKXKWKVKUNNNNNNNNNNNNNNNKCKBKAK@K?K@KAKBNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKkKjKiKhKgKfKeNNNNNNNNNNNNNNKTKSKRKQKPKOKNKMKLKKKJKIKHKGKFKEKDKCKBKAK@KAKBKCNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKlKkKjKiKhKgKfNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKEKDKCKBKAKBKCKDNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKmKlKkKjKiKhKgNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKEKDKCKBKCKDKENNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKnKmKlKkKjKiKhNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKFKEKDKCKDKEKFNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKoKnKmKlKkKjKiNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKGKFKEKDKEKFKGNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKpKoKnKmKlKkKjNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKIKHKGKFKEKFKGKHNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKqKpKoKnKmKlKkNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKJKIKHKGKFKGKHKINNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKJKIKHKGKHKIKJNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�Tiles�}�(K }�(K �Tile�jB/  ��)��}�(j,,  j]-  j&,  ]�j0,  K j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�K%aj0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLub�      KMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�K&aj0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�K'aj0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�K(aj0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�K)aj0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK	}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K	j1,  KOubuK
}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K
j1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�K*aj0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;�      jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�K+aj0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�K,aj0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�K-aj0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�K.aj0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�K/aj0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�K0aj0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�K1aj0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�K2aj0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�K3aj0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�K4aj0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  Kj1,  KOubuK }�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K j1,  KOubuK!}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K!j1,  KOubuK"}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K"j1,  KOubuK#}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K#j1,  KOubuK$}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K$j1,  KOubuK%}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K%j1,  KOubuK&}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�K5aj0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K&j1,  KOubuK'}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  �      K'j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K'j1,  KOubuK(}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K(j1,  KOubuK)}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K)j1,  KOubuK*}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K*j1,  KOubuK+}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K+j1,  KOubuK,}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K,j1,  KOubuK-}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K-j1,  KOubuK.}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K.j1,  KOubuK/}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�K6aj0,  K/j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K/j1,  KOubuK0}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�K8aj0,  K0j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K0j1,  KOubuK1}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K1j1,  KOubuK2}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K2j1,  KOubuK3}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K3j1,  KOubuK4}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�K9aj0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K4j1,  KOubuK5}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�K:aj0,  K5j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�K;aj0,  K5j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�K<aj0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�K=aj0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K5j1,  KOubuK6}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�K>aj0,  K6j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K6j1,  KOubuK7}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K7j1,  KOubuK8}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K8j1,  KOubuK9}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  �      ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K9j1,  KOubuK:}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K:j1,  KOubuK;}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K;j1,  KOubuK<}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K<j1,  KOubuK=}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�K?aj0,  K=j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K=j1,  KOubuK>}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�K@aj0,  K>j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K>j1,  KOubuK?}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�KCaj0,  K?j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K?j1,  KOubuK@}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�KDaj0,  K@j1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  K@j1,  KOubuKA}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�KEaj0,  KAj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KAj1,  KOubuKB}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�KFaj0,  KBj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KBj1,  KOubuKC}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�KGaj0,  KCj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KCj1,  KOubuKD}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�KHaj0,  KDj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KDj1,  KOubuKE}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�K7aj0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KEj1,  KOubuKF}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KFj1,  KOubuKG}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KGj1,  KOubuKH}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KHj1,  KOubuKI}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KIj1,  KOubuKJ}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KJj1,  KOubuKK}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  �      j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KKj1,  KOubuKL}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KLj1,  KOubuKM}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KMj1,  KOubuKN}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KNj1,  KOubuKO}�(K jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubK	jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K	ubK
jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K
ubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KubK jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K ubK!jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K!ubK"jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K"ubK#jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K#ubK$jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K$ubK%jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K%ubK&jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K&ubK'jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K'ubK(jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K(ubK)jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K)ubK*jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K*ubK+jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K+ubK,jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K,ubK-jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K-ubK.jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K.ubK/jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K/ubK0jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K0ubK1jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K1ubK2jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K2ubK3jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K3ubK4jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K4ubK5jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K5ubK6jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K6ubK7jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K7ubK8jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K8ubK9jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K9ubK:jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K:ubK;jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K;ubK<jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K<ubK=jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K=ubK>jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K>ubK?jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K?ubK@jC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  K@ubKAjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KAubKBjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KBubKCjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KCubKDjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KDubKEjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KEubKFjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KFubKGjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KGubKHjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KHubKIjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KIubKJjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KJubKKjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KKubKLjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KLubKMjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KMubKNjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KNubKOjC/  )��}�(j,,  j]-  j&,  ]�j0,  KOj1,  KOubuu�	enemyList�]�(j�,  j�,  e�master_Changed_Tiles�]�(]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KDKe]�(KEKe]�(KDKe]�(KEKe]�(KDKe]�(KEKe]�(KDKe]�(KEKe]�(KDKe]�(KEKe]�(KDKe]�(KEKe]�(KDKe]�(KEKe]�(KEKe]�(KDKe]�(KEKe]�(KEKe]�(KDKe]�(KEKe]�(KEKe]�(KEKe]�(KDKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KDKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KDKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEK
e]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KFKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KEKe]�(KFKe]�(KEKe]�(KEKe]�(KFKe]�(KEKe]�(KEKe]�(KEKe]�(KFKe]�(KEKe]�(KFKe]�(KEKe]�(KEKe]�(KFKe]�(KEKe]�(KFKe]�(KEKe]�(KFKe]�(KEKe]�(KFKe]�(KEKe]�(KFKe]�(KFKe]�(KEKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKe]�(KDKe]�(KFKeej9,  j[-  �djikstra_Player�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�P�     G�P�     G�P      G�P�     G�P�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�P�     G�P      G�O�     G�P      G�P�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�P      G�O�     G�N�     G�O�     G�P      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�O�     G�N�     G�N      G�N�     G�O�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�N�     G�N      G�M@     G�N      G�N�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�N      G�M@     G�L�     G�M@     G�N      G�N�     G�O�     G�P      G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      G�S�     G�S�     G�T@     NNNNNNNNNNNNG�U`     G�U      G�T�     G�T@     G�S�     G�T@     G�T�     G�U      G�U`     G�U�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�M@     G�L�     G�K�     G�L�     G�M@     NNNNNNNNNNNNNG�T�     NNNNNNNNNNNNG�U      G�T�     G�T@     G�S�     G�S�     G�S�     G�T@     G�T�     G�U      G�U`     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNG�L�     G�K�     G�K      G�K�     G�L�     NNNNNNNNNNNNNG�U      NNNNNNNNNNNNNNNNG�S      G�S�     G�S�     G�T@     G�T�     G�U      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�J@     G�K      G�K�     NNNNNNNNNNNNNG�U`     NNNNNNNNNNNNNNNNG�R�     G�S      G�S�     G�S�     G�T@     G�T�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�I�     G�J@     G�K      NNNNNNNNNNNNNG�U�     NNNNNNNNNNNNNNNNG�R`     G�R�     G�S      G�S�     G�S�     G�T@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�H�     NNNNNNNNNNNNNNNG�V      NNNNNNNNNNNNNG�Q�     NNG�R      G�R`     G�R�     G�S      G�S�     G�S�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�H      NNNNNNNNNNNNNNNK NNNNNNNNNNNNG�Q�     G�Q@     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      G�S�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�G@     NNNNNNNNNNNNNNNG�V      NNNNNNNNNNNNG�Q@     G�P�     G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     G�S      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�F�     NNNNNNNNNNNNNNNG�U�     G�U`     G�U      G�T�     G�T@     G�S�     G�S�     G�S      G�R�     G�R`     G�R      G�Q�     G�Q@     G�P�     G�P�     G�P      G�P�     G�P�     G�Q@     G�Q�     G�R      G�R`     G�R�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNG�E�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�O�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�B�     G�C�     G�D@     G�E      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�N�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�B      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�N      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�A@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�M@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�@�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�L�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�?�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�K�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�>      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�K      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�<�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�J@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�;      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�I�     G�J@     G�K      G�K�     G�L�     G�M@     G�N      G�N�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�>      G�<�     G�;      G�9�     G�8      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�H�     G�I�     G�J@     G�K      G�K�     G�L�     G�M@     G�N      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�<�     G�;      G�9�     G�8      G�6�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�H      G�H�     G�I�     G�J@     G�K      G�K�     G�L�     G�M@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�;      G�9�     G�8      G�6�     G�5      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�G@     G�H      G�H�     G�I�     G�J@     G�K      G�K�     G�L�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�9�     G�8      G�6�     G�5      G�3�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�F�     G�G@     G�H      G�H�     G�I�     G�J@     G�K      G�K�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�8      G�6�     G�5      G�3�     G�2      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�E�     G�F�     G�G@     G�H      G�H�     G�I�     G�J@     G�K      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�6�     G�5      G�3�     G�2      G�0�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�E      G�E�     G�F�     G�G@     G�H      G�H�     G�I�     G�J@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�5      G�3�     G�2      G�0�     G�.      NNNNNNNNNNNNNNNG�.      G�0�     G�2      G�3�     G�5      G�6�     G�8      G�9�     G�;      G�<�     G�>      G�?�     G�@�     G�A@     G�B      G�B�     G�C�     G�D@     G�E      G�E�     G�F�     G�G@     G�H      G�H�     G�I�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNG�0�     G�.      G�+      NNNNNNNNNNNNNNNG�+      NNNNNNNNNNNNNNNNNG�E�     G�F�     G�G@     G�H      G�H�     G�I�     G�J@     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNG�.      G�+      G�(      G�%      G�"      G�      G�      G�      G�      G��      G�       G��      G�      G�      G�      G�      G�"      G�%      G�(      NNNNNNNNNNNNNNNNNNG�G@     G�H      G�H�     G�I�     G�J@     G�K      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�	decorList�]�(j4,  j�-  jA.  e�	textSpace��Ornate mosaic floor
��SeenMap�]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K ee�maze�]�(]�(�#�j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  �.�j�{  j�-  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j.,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j,  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�-  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j.,  j.,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j.,  j.,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  jF,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j.,  j.,  j�{  j�{  j�{  j�-  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j.,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j<,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j<,  j<,  j<,  j<,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j<,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  �      j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  jF,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  jq,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  jV,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  jV,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j.,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  ee�levelManager�j�+  �	thePlayer�j�,  �consumeList�]�(j�+  j�+  j�+  j�+  j�+  e�	tilesSeen�]��
stairsDown�]�(KKe�djikstra_Stairs_Up�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK6K5K4K3K2NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK5K4K3K2K1NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK4K3K2K1K0NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK3K2K1K0K/NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK2K1K0K/K.NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK1K0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KNNNNNNNNNNNNK
K	KKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK2K1K0K/K.NNNNNNNNNNNNNKNNNNNNNNNNNNK	KKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK3K2K1K0K/NNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK2K1K0NNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK3K2K1NNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKKK KKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK4NNNNNNNNNNNNNNNKNNNNNNNNNNNNNKNNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK5NNNNNNNNNNNNNNNKNNNNNNNNNNNNKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK6NNNNNNNNNNNNNNNKNNNNNNNNNNNNK	KKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK7NNNNNNNNNNNNNNNKKKKKKKKKKKKKK
K	KKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK8NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK	NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK<K;K:K9NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK
NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK=NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK?NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK@NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKANNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKBNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKGKFKEKDKCNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKFKEKDKCKBNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKEKDKCKBKANNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKDKCKBKAK@NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKCKBKAK@K?NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKBKAK@K?K>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKAK@K?K>K=NNNNNNNNNNNNNNNK)K(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNK>K=K<NNNNNNNNNNNNNNNK*NNNNNNNNNNNNNNNNNKKKKKKK NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNK=K<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+NNNNNNNNNNNNNNNNNNKKKKK K!NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�	gameState�h�djikstra_Player_Adj�]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK5K4K3K2K1NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK4K3K2K1K0NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK3K2K1K0K/NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK2K1K0K/K.NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK1K0K/K.K-NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK0K/K.K-K,K+K*K)K(K'K&K%K$K#K"K!K KKNNNNNNNNNNNNK	KKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK1K0K/K.K-NNNNNNNNNNNNNKNNNNNNNNNNNNKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNK2K1K0K/K.NNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK1K0K/NNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKKK KKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK2K1K0NNNNNNNNNNNNNKNNNNNNNNNNNNNNNNKK KK KKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK3NNNNNNNNNNNNNNNKNNNNNNNNNNNNNKNNKKK KKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK4NNNNNNNNNNNNNNNKNNNNNNNNNNNNKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK5NNNNNNNNNNNNNNNKNNNNNNNNNNNNKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK6NNNNNNNNNNNNNNNKKKKKKKKKKKKK
K	KKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNK7NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK;K:K9K8NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK	NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK<NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNK
NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK=NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK?NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNK@NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKANNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKBNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKFKEKDKCKBNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKEKDKCKBKANNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKDKCKBKAK@NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKCKBKAK@K?NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKBKAK@K?K>NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKAK@K?K>K=NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK@K?K>K=K<NNNNNNNNNNNNNNNK(K'K&K%K$K#K"K!K KKKKKKKKKKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNK=K<K;NNNNNNNNNNNNNNNK)NNNNNNNNNNNNNNNNNKKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNK<K;K:K9K8K7K6K5K4K3K2K1K0K/K.K-K,K+K*NNNNNNNNNNNNNNNNNNKKKKKK NNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNee�djikstra_Player_Away�j:{  j7,  �2B: Dark Crypt��
messageSys��
MessageSys��Messages���)��}�(�messages�]�(�Kyle acquired 19 coins��Kyle picked up Green Herb��'Kyle picked up Scroll of Lightning Bolt��Kyle picked up +1 Iron Helm��Kyle picked up Bomb��Kyle picked up Longsword��Kyle picked up Longsword��Kyle picked up +1 Leather Helm��Zombie dropped Longsword��Zombie dropped +1 Leather Helm��Zombie was killed by Kyle��Zombie is afraid!��Kyle attacked Zombie for 3��Zombie attacked Kyle for 5��Kyle attacked Zombie for 3��Zombie attacked Kyle for 5��Kyle picked up +1 Iron Helm��Zombie attacked Kyle for 5��Skeleton Knight dropped Bomb��!Skeleton Knight dropped Longsword��$Skeleton Knight dropped +1 Iron Helm��"Skeleton Knight was killed by Kyle��Skeleton Knight is afraid!��#Kyle attacked Skeleton Knight for 2��#Skeleton Knight attacked Kyle for 6��Kyle missed Skeleton Knight��#Skeleton Knight attacked Kyle for 6��#Kyle attacked Skeleton Knight for 2��#Skeleton Knight attacked Kyle for 6��#Kyle attacked Skeleton Knight for 2��Skeleton Knight missed Kyle��#Kyle attacked Skeleton Knight for 2��#Skeleton Knight attacked Kyle for 6��Kyle acquired 13 coins��Kyle picked up Longsword��Kyle picked up Chain Shirt��Kyle acquired 6 Arrows��Kyle acquired 9 coins��Kyle picked up Green Herb��Kyle picked up Iron Helm��Kyle picked up Buckler��Kyle picked up Bomb��Kyle acquired 4 coins��Kyle picked up Longsword��Kyle picked up Longsword��Kyle picked up Iron Helm��Skeleton Knight dropped Bomb��!Skeleton Knight dropped Longsword��!Skeleton Knight dropped Iron Helm��"Skeleton Knight was killed by Kyle��Skeleton Knight is afraid!��#Kyle attacked Skeleton Knight for 3��#Skeleton Knight attacked Kyle for 4��#Kyle attacked Skeleton Knight for 3��#Skeleton Knight attacked Kyle for 4��Kyle picked up Iron Helm��#Skeleton Knight attacked Kyle for 4��"Skeleton Knight dropped Gold Coins��!Skeleton Knight dropped Longsword��!Skeleton Knight dropped Iron Helm��"Skeleton Knight was killed by Kyle��Skeleton Knight is afraid!��#Kyle attacked Skeleton Knight for 3��#Skeleton Knight attacked Kyle for 4��#Kyle attacked Skeleton Knight for 3��Kyle waited...��Kyle acquired 7 coins��Kyle picked up Longsword��Kyle picked up Iron Helm��"Skeleton Knight dropped Gold Coins��!Skeleton Knight dropped Longsword��!Skeleton Knight dropped Iron Helm��"Skeleton Knight was killed by Kyle��Skeleton Knight is afraid!��#Kyle attacked Skeleton Knight for 3��#Skeleton Knight attacked Kyle for 4��#Kyle attacked Skeleton Knight for 3��#Skeleton Knight attacked Kyle for 4��Kyle picked up Green Herb��'Kyle picked up Scroll of Lightning Bolt��Kyle picked up Longsword��Kyle picked up Longsword��Kyle picked up Iron Helm��0Skeleton Knight dropped Scroll of Lightning Bolt��!Skeleton Knight dropped Longsword��!Skeleton Knight dropped Iron Helm��"Skeleton Knight was killed by Kyle��Skeleton Knight is afraid!��#Kyle attacked Skeleton Knight for 3��#Skeleton Knight attacked Kyle for 4��#Kyle attacked Skeleton Knight for 3��Kyle acquired 15 coins��Kyle picked up Iron Helm��Kyle picked up Wooden Shield��Kyle picked up Iron Helm��Kyle picked up Leather Helm��Zombie dropped Longsword��Zombie dropped Leather Helm��Zombie was killed by Kyle��Zombie is afraid!��Kyle attacked Zombie for 3��Zombie attacked Kyle for 3��Kyle attacked Zombie for 3��Zombie attacked Kyle for 3��Player Ready: Kyle��
Game Start�e�messageLimit�M��retrieveLimit�Kub�SeesMap�]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K KK K KKKKKKKKK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K KKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K KK K KKKKKKKKK K KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K ee�inSeed�M��textWall��Ornate stone wall
�ubj-,  j�,  j/,  K7j0,  KEj1,  Kj(,  j�,  j7,  j�,  ub�skillPoints�Kj�,  ]�j�,  Kj�,  KdjB,  ]�(KKYK�ej7,  �Kyle�ubj7,  j�,  ubKj),  )��}�(j,,  j�+  j-,  j.,  j/,  Kj0,  Kj1,  Kj(,  jA.  )��}�(j7,  jD.  j9,  j�}  j-,  j.,  ubj7,  jD.  ubK	j�,  K
j),  )��}�(j,,  j�+  j-,  j,  j/,  K
j0,  Kj1,  Kj(,  j�,  )��}�(jd,  Kj�,  K j-,  j,  j�,  K(j�,  ]�(j�}  j),  )��}�(j,,  j�+  j-,  j,  j/,  Kj0,  Kj1,  K"j(,  j�,  )��}�(jd,  Kj�,  K j-,  j,  j�,  K(j�,  ]�(j�}  j�}  ej�,  Kj�,  �j�,  j,  )��}�(jn,  K
jd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  j�,  ubj�,  K j�,  Kj�,  K j�,  K j�,  K	j�,  Kj�,  Kj�,  Nj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  js,  ubj�,  Kj�,  �j�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  Kjr,  �j7,  j ,  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  j�}  j�,  Kdj�,  ]�j�,  K jB,  j�,  j7,  j�,  ubj7,  j�,  ubej�,  Kj�,  �j�,  j,  )��}�(jn,  K
jd,  KjI,  �jJ,  �jo,  KjL,  j�,  jB,  jM,  j-,  jq,  jr,  �j7,  j�,  ubj�,  K j�,  Kj�,  K j�,  K j�,  K	j�,  Kj�,  Kj�,  Nj�,  G        j�,  �j�,  �j[,  ]�jp,  j,  )��}�(jn,  Kjd,  KjI,  �jJ,  �jo,  KjL,  jp,  jB,  jM,  j-,  jq,  jr,  �j7,  js,  ubj�,  Kj�,  �j�,  Nj�,  K j�,  Nj�,  j,  )��}�(jd,  Kj-,  jq,  jL,  j�,  jI,  �jJ,  �j�,  �j�,  Kj�,  Kjo,  Kj�,  Kj�,  �jB,  jM,  j�,  Kjr,  �j7,  j ,  ubj�,  Njn,  K j�,  �j�,  �j�,  K j�,  Nj�,  Kj�,  Kj�,  Nj�,  �j�,  ]�j9,  j�}  j�,  Kdj�,  ]�j�,  K jB,  j�,  j7,  j�,  ubj7,  j�,  ubKj�}  Kj),  )��}�(j,,  j�+  j-,  jV,  j/,  Kj0,  Kj1,  K	j(,  jX,  )��}�(j[,  ]�j9,  j�}  jB,  jM,  j-,  jV,  j7,  jW,  ubj7,  jW,  ubKj),  )��}�(j,,  j�+  j-,  jF,  j/,  Kj0,  K!j1,  Kj(,  j-  j7,  jO,  ubKj),  )��}�(j,,  j�+  j-,  j.,  j/,  Kj0,  K(j1,  K%j(,  j4,  )��}�(j7,  j8,  j9,  j�}  j-,  j.,  ubj7,  j8,  ubKj),  )��}�(j,,  j�+  j-,  j�-  j/,  Kj0,  K(j1,  K)j(,  j�-  )��}�(j,,  j�+  j9,  j�}  j/,  J����j0,  K(j�,  Kj(,  Nj1,  K)j7,  j�,  ubj7,  j�-  ubKj),  )��}�(j,,  j�+  j-,  jV,  j/,  Kj0,  K)j1,  K'j(,  jX,  )��}�(j[,  ]�j9,  j�}  jB,  jM,  j-,  jV,  j7,  jW,  ubj7,  jW,  ubKj),  )��}�(j,,  j�+  j-,  jV,  j/,  Kj0,  K-j1,  K%j(,  jX,  )��}�(j[,  ]�j9,  j�}  jB,  jM,  j-,  jV,  j7,  jW,  ubj7,  jW,  ubKj),  )��}�(j,,  j�+  j-,  jq,  j/,  Kj0,  Kj1,  K	j(,  j-  j7,  j�,  ubKj),  )��}�(j,,  j�+  j-,  jq,  j/,  Kj0,  Kj1,  K	j(,  j-  j7,  j ,  ubKj),  )��}�(j,,  j�+  j-,  jq,  j/,  Kj0,  Kj1,  Kj(,  j-  j7,  j�,  ubKj),  )��}�(j,,  j�+  j-,  jq,  j/,  Kj0,  Kj1,  Kj(,  j-  j7,  j ,  ubKj),  )��}�(j,,  j�+  j-,  jj,  j/,  Kj0,  Kj1,  Kj(,  j-  j7,  j-  ubKj),  )��}�(j,,  j�+  j-,  jq,  j/,  Kj0,  K*j1,  Kj(,  j-  j7,  j�,  ubKj),  )��}�(j,,  j�+  j-,  jq,  j/,  Kj0,  K*j1,  Kj(,  j-  j7,  j ,  ubKj),  )��}�(j,,  j�+  j-,  jy,  j/,  Kj0,  K*j1,  Kj(,  ju,  )��}�(jI,  �jJ,  �j9,  NjL,  jJ,  jB,  jx,  j-,  jy,  jz,  Kj7,  j{,  ubj7,  j{,  ubKj),  )��}�(j,,  j�+  j-,  jq,  j/,  Kj0,  K,j1,  K$j(,  j-  j7,  j�,  ubK j),  )��}�(j,,  j�+  j-,  jq,  j/,  K j0,  K,j1,  K$j(,  j!-  j7,  j ,  ubK!j),  )��}�(j,,  j�+  j-,  jy,  j/,  K!j0,  K,j1,  K$j(,  ju,  )��}�(jI,  �jJ,  �j9,  NjL,  jJ,  jB,  jx,  j-,  jy,  jz,  Kj7,  j{,  ubj7,  j{,  ubK"j),  )��}�(j,,  j�+  j-,  jq,  j/,  K"j0,  K+j1,  K$j(,  j-  j7,  j�,  ubK#j),  )��}�(j,,  j�+  j-,  jq,  j/,  K#j0,  K+j1,  K$j(,  j#-  j7,  j ,  ubK$j),  )��}�(j,,  j�+  j-,  j'-  j/,  K$j0,  K+j1,  K$j(,  j%-  j7,  j)-  ubuj�.  ]�(]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKK K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKKK K K K K KKKKKKKKKKKK KKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKKKKKKKKKK KKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKKKKKKKKKK KKKKKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKKKKKKKKKK KKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K K K K K K K K K K K K K KKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKK K K K KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKK K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKK KKKKKKKKKKKKKK KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKK KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKK KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKK KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K K K K K K K K K K K K KKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKKKKKKKKK K K K K K K KKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKK K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K KKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKK K K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K KKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKe]�(KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKeej�.  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNK[KZKYKZNNNNNNNNNNNKfKgKhKiKjKkKlKmKnKoKpKqKpKoKnKoKpKqKrNNNNNNNNNNNNNNNNNNNNNNe]�(NNNK[KZKYKXKYNNNNNNNNNNNKeNNNNNNNNNNKpKoKnKmKnKoKpKqNNNNNNNNNNNNNNNNNNNNNNe]�(NNK[KZKYKXKWKXNNNNNNNNNNNKdNNNNNNNNNNKoKnKmKlKmKnKoKpNNNNNNNNNNNNNNNNNNNNNNe]�(NNKZKYKXKWKVKWNNNNNNNNNNNKcNNNNNNNNNNKnKmKlKkKlKmKnKoNNNNNNNNNNNNNNNNNNNNNNe]�(NNKYKXKWKVKUKVNNNNNNNNNNNKbNNNNNNNNNNNKlKkKjKkKlKmKnNNNNNNNNNNNNNNNNNNNNNNe]�(NNKXKWKVKUKTKUKVKWKXKYKZK[K\K]K^K_K`KaNNNNNNNNNNNNKjKiKjKkKlKmNNNNNNNNNNNNNNNNNNNNNNe]�(NNKWKVKUKTKSKTNNNNNNNNNNNNNNNNNNNNNNNNNKhNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKVKUKTKSKRKSNNNNNNNNNNNNNNNNNNNNNNNNNKgNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKUKTKSKRKQKRNNNNNNNNNNNNNNNNNNNNNNNNNKfNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKPNNNNNNNNNNNNNNNNNNNNNNNNNNKeNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKONNNNNNNNNNNNNNNNNNNNNNNNNNKdNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNKcNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKMNNNNNNNNNNNNNNNNNNNNNNNNNNKbNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKLNNNNNNNNNNNNNNNNNNNNNNNNNNKaNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKKKJKIKHNNNNNNNNNNNNNNNNNNNNNNNK`NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKGNNNNNNNNNNNNNNNNNNNNNNNK_NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKFNNNNNNNNNNNNNNNNNNNNNNNK^NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKENNNNNNNNNNNNNNNNNNNNNNNK]NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKDNNNNNNNNNNNNNNNNNNNNNNNK\NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKCNNNNNNNNNNNNNNNNNNNNNNNK[NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKBNNNNNNNNNNNNNKPKQKRKSKTKUKVKWKXKYKZK[K\K]NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKANNNNNNNNNNNNNKONNNNNNKXKYKZK[K\K]K^NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK>K?K@KAKBKCNNNNNNNNNNKNNNNNNNKYKZK[K\K]K^K_NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK=K>K?K@KAKBNNNNNNNNNNKMNNNNNNKZK[K\K]K^K_K`NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK<K=K>K?K@KANNNNNNNNNNKLNNNNNNK[K\K]K^K_K`KaNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK;K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKNNNNNNK\K]K^K_K`KaKbNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK:K;K<K=K>K?NNNNNNNNNNNNNNNNNK]K^K_K`KaKbKcNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK9K:K;K<K=K>NNNNNNNNNNNNNNNNNK^K_K`KaKbKcKdNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK8K9K:K;K<K=NNNNNNNNNNNNNNNNNK_K`KaKbKcKdKeNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK7K8K9K:K;K<NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK6NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK5NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK4NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK3NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNK.K/K0K1NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK-NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKK NNNNNNNNNNNNNNNNNNe]�(NNNNK,NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK+K*K)K(K'NNNNNNNNNNNNNNNNNNNNNNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK*K)K(K'K&K%K$K#K"K!K KKKKKNNNNNNNNNNNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK+K*K)K(K'NNNNNNNNNNKKKKKKKKKKKKKKKKK
K	KKKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK,K+K*K)K(NNNNNNNNNNNNNNNNNNNNNNNNNNNK
K	KKKKNNNNNNNNNNNNNNNNNNe]�(NNNNK-K,K+K*K)NNNNNNNNNNNNNNNNNNNNNNNNNNNKK
K	KKKNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKKK
K	KKNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej?/  }�(K }�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  �      ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�K aj0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�Kaj0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�Kaj0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�Kaj0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�Kaj0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�Kaj0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�Kaj0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�Kaj0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�K	aj0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK	}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K	j1,  K;ubuK
}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K
j1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�K
aj0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�Kaj0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  �      j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�Kaj0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  Kj1,  K;ubuK }�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K j1,  K;ubuK!}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K!j1,  K;ubuK"}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K"j1,  K;ubuK#}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K#j1,  K;ubuK$}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K$j1,  K;ubuK%}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K%j1,  K;ubuK&}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K&j1,  K;ubuK'}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K'j1,  K;ubuK(}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�Kaj0,  K(j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�(KKej0,  K(j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K(j1,  K;ubuK)}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�Kaj0,  K)j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K)j1,  K;ubuK*}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K*j1,  K;ubuK+}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K+j1,  K;ubuK,}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K,j1,  K;ubuK-}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�Kaj0,  K-j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K-j1,  K;ubuK.}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K.j1,  K;ubuK/}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K/j1,  K;ubuK0}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K0j1,  K;ubuK1}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K1j1,  K;ubuK2}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K2j1,  K;ubuK3}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  �       K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K3j1,  K;ubuK4}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K4j1,  K;ubuK5}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K5j1,  K;ubuK6}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K6j1,  K;ubuK7}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K7j1,  K;ubuK8}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K8j1,  K;ubuK9}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K9j1,  K;ubuK:}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K:j1,  K;ubuK;}�(K jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubK	jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K	ubK
jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K
ubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubKjC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  KubK jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K ubK!jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K!ubK"jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K"ubK#jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K#ubK$jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K$ubK%jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K%ubK&jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K&ubK'jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K'ubK(jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K(ubK)jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K)ubK*jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K*ubK+jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K+ubK,jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K,ubK-jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K-ubK.jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K.ubK/jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K/ubK0jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K0ubK1jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K1ubK2jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K2ubK3jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K3ubK4jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K4ubK5jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K5ubK6jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K6ubK7jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K7ubK8jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K8ubK9jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K9ubK:jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K:ubK;jC/  )��}�(j,,  j�+  j&,  ]�j0,  K;j1,  K;ubuuj�z  j�z  j�z  ]�(]�(K'K'e]�(K&K&e]�(K'K)e]�(K&K*e]�(K'K'e]�(K&K&e]�(K'K)e]�(K&K*e]�(K'K'e]�(K&K&e]�(K'K)e]�(K&K*e]�(K'K'e]�(K&K&e]�(K'K)e]�(K'K*e]�(K'K'e]�(K'K&e]�(K&K%e]�(K'K)e]�(K'K*e]�(K'K'e]�(K'K&e]�(K&K%e]�(K'K)e]�(K'K*e]�(K'K'e]�(K'K&e]�(K&K%e]�(K(K)e]�(K'K*e]�(K(K'e]�(K'K&e]�(K'K%e]�(K(K)e]�(K'K*e]�(K(K'e]�(K'K&e]�(K'K%e]�(K(K)e]�(K'K*e]�(K(K'e]�(K'K&e]�(K'K%e]�(K(K)e]�(K(K*e]�(K(K'e]�(K(K&e]�(K'K%e]�(K(K)e]�(K(K*e]�(K(K'e]�(K(K&e]�(K(K%e]�(K(K$e]�(K(K)e]�(K(K*e]�(K(K'e]�(K(K&e]�(K(K%e]�(K(K$e]�(K(K)e]�(K(K*e]�(K(K'e]�(K(K&e]�(K(K%e]�(K(K$e]�(K(K)e]�(K(K*e]�(K(K'e]�(K(K&e]�(K)K%e]�(K)K$e]�(K)K#e]�(K(K)e]�(K(K*e]�(K(K'e]�(K)K&e]�(K)K%e]�(K)K$e]�(K)K#e]�(K(K)e]�(K(K*e]�(K(K'e]�(K)K&e]�(K)K%e]�(K)K$e]�(K*K#e]�(K(K)e]�(K)K*e]�(K(K'e]�(K)K&e]�(K)K%e]�(K*K$e]�(K*K#e]�(K(K)e]�(K)K*e]�(K)K'e]�(K)K&e]�(K*K%e]�(K*K$e]�(K+K#e]�(K(K)e]�(K)K*e]�(K)K'e]�(K)K&e]�(K*K%e]�(K*K$e]�(K+K#e]�(K)K)e]�(K)K*e]�(K)K'e]�(K)K&e]�(K*K%e]�(K+K$e]�(K+K#e]�(K)K)e]�(K)K*e]�(K)K'e]�(K*K&e]�(K*K%e]�(K+K$e]�(K,K#e]�(K-K"e]�(K)K)e]�(K)K*e]�(K)K'e]�(K*K&e]�(K+K%e]�(K+K$e]�(K,K#e]�(K-K"e]�(K)K)e]�(K*K*e]�(K)K'e]�(K*K&e]�(K+K%e]�(K,K$e]�(K-K#e]�(K)K)e]�(K*K*e]�(K)K'e]�(K*K&e]�(K+K%e]�(K,K$e]�(K-K#e]�(K)K)e]�(K*K*e]�(K'K'e]�(K&K&e]�(K)K'e]�(K*K&e]�(K+K%e]�(K,K$e]�(K-K#e]�(K'K'e]�(K&K&e]�(K)K'e]�(K*K&e]�(K+K%e]�(K,K$e]�(K-K#e]�(K'K'e]�(K&K&e]�(K)K'e]�(K*K&e]�(K+K&e]�(K,K%e]�(K-K$e]�(K.K#e]�(K'K'e]�(K&K&e]�(K)K'e]�(K*K'e]�(K+K&e]�(K,K%e]�(K-K$e]�(K.K$e]�(K/K#e]�(K'K'e]�(K&K'e]�(K)K'e]�(K*K'e]�(K+K&e]�(K,K%e]�(K-K%e]�(K.K$e]�(K/K#e]�(K'K'e]�(K&K'e]�(K)K'e]�(K*K'e]�(K+K&e]�(K,K&e]�(K-K%e]�(K.K%e]�(K/K$e]�(K0K#e]�(K'K'e]�(K&K'e]�(K)K(e]�(K*K'e]�(K+K'e]�(K,K&e]�(K-K&e]�(K.K%e]�(K/K%e]�(K0K$e]�(K'K(e]�(K&K'e]�(K)K(e]�(K*K'e]�(K+K'e]�(K,K&e]�(K-K&e]�(K.K&e]�(K/K%e]�(K0K%e]�(K'K(e]�(K&K'e]�(K)K(e]�(K*K'e]�(K+K'e]�(K,K'e]�(K-K&e]�(K.K&e]�(K/K&e]�(K0K%e]�(K'K(e]�(K&K'e]�(K)K(e]�(K*K(e]�(K+K'e]�(K,K'e]�(K-K'e]�(K.K'e]�(K/K&e]�(K0K&e]�(K'K(e]�(K&K(e]�(K)K(e]�(K*K(e]�(K+K(e]�(K,K'e]�(K-K'e]�(K.K'e]�(K/K'e]�(K0K'e]�(K'K(e]�(K&K(e]�(K)K(e]�(K*K(e]�(K+K(e]�(K,K(e]�(K-K(e]�(K.K(e]�(K/K'e]�(K0K'e]�(K'K(e]�(K&K(e]�(K)K(e]�(K*K(e]�(K+K(e]�(K,K(e]�(K-K(e]�(K.K(e]�(K/K(e]�(K0K(e]�(K'K(e]�(K&K(e]�(K)K(e]�(K*K(e]�(K+K(e]�(K,K(e]�(K-K(e]�(K.K(e]�(K/K)e]�(K0K)e]�(K'K(e]�(K&K(e]�(K)K(e]�(K*K(e]�(K+K(e]�(K,K)e]�(K-K)e]�(K.K)e]�(K/K)e]�(K0K)e]�(K'K(e]�(K&K)e]�(K)K(e]�(K*K(e]�(K+K)e]�(K,K)e]�(K-K)e]�(K.K)e]�(K/K*e]�(K'K(e]�(K&K)e]�(K)K(e]�(K*K)e]�(K+K)e]�(K,K)e]�(K-K*e]�(K'K(e]�(K&K)e]�(K)K(e]�(K*K)e]�(K+K)e]�(K,K*e]�(K'K)e]�(K&K)e]�(K)K(e]�(K*K)e]�(K+K)e]�(K,K*e]�(K'K)e]�(K&K)e]�(K)K)e]�(K*K)e]�(K+K*e]�(K'K)e]�(K&K)e]�(K)K)e]�(K*K)e]�(K+K*e]�(K'K)e]�(K&K*e]�(K)K)e]�(K*K)e]�(K+K*e]�(K'K)e]�(K&K*e]�(K)K)e]�(K*K*e]�(K'K)e]�(K&K*e]�(K)K)e]�(K*K*e]�(K'K)e]�(K&K*e]�(K)K)e]�(K*K*e]�(K(K(e]�(K(K)eej9,  j�,  j9{  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNG�`�     G�`�     G�`�     G�`�     NNNNNNNNNNNG�b�     G�c      G�cP     G�c�     G�c�     G�c�     G�d     G�d@     G�dp     G�d�     G�d�     G�e      G�d�     G�d�     G�dp     G�d�     G�d�     G�e      K NNNNNNNNNNNNNNNNNNNNNNe]�(NNNG�`�     G�`�     G�`�     G�`P     G�`�     NNNNNNNNNNNG�b�     NNNNNNNNNNG�d�     G�d�     G�dp     G�d@     G�dp     G�d�     G�d�     G�e      NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`�     G�`�     G�`P     G�`      G�`P     NNNNNNNNNNNG�b�     NNNNNNNNNNG�d�     G�dp     G�d@     G�d     G�d@     G�dp     G�d�     G�d�     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`�     G�`P     G�`      G�_�     G�`      NNNNNNNNNNNG�b`     NNNNNNNNNNG�dp     G�d@     G�d     G�c�     G�d     G�d@     G�dp     G�d�     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`�     G�`P     G�`      G�_�     G�_�     G�_�     NNNNNNNNNNNG�b0     NNNNNNNNNNNG�d     G�c�     G�c�     G�c�     G�d     G�d@     G�dp     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`P     G�`      G�_�     G�_�     G�_      G�_�     G�_�     G�`      G�`P     G�`�     G�`�     G�`�     G�a     G�a@     G�ap     G�a�     G�a�     G�b      NNNNNNNNNNNNG�c�     G�c�     G�c�     G�c�     G�d     G�d@     NNNNNNNNNNNNNNNNNNNNNNe]�(NNG�`      G�_�     G�_�     G�_      G�^�     G�_      NNNNNNNNNNNNNNNNNNNNNNNNNG�cP     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�_�     G�_�     G�_      G�^�     G�^`     G�^�     NNNNNNNNNNNNNNNNNNNNNNNNNG�c      NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNG�_�     G�_      G�^�     G�^`     G�^      G�^`     NNNNNNNNNNNNNNNNNNNNNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�]�     NNNNNNNNNNNNNNNNNNNNNNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�]@     NNNNNNNNNNNNNNNNNNNNNNNNNNG�b�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�\�     NNNNNNNNNNNNNNNNNNNNNNNNNNG�b`     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�\�     NNNNNNNNNNNNNNNNNNNNNNNNNNG�b0     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�\      NNNNNNNNNNNNNNNNNNNNNNNNNNG�b      NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNG�[�     G�[`     G�[      G�Z�     NNNNNNNNNNNNNNNNNNNNNNNG�a�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�Z@     NNNNNNNNNNNNNNNNNNNNNNNG�a�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�Y�     NNNNNNNNNNNNNNNNNNNNNNNG�ap     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�Y�     NNNNNNNNNNNNNNNNNNNNNNNG�a@     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�Y      NNNNNNNNNNNNNNNNNNNNNNNG�a     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�X�     NNNNNNNNNNNNNNNNNNNNNNNG�`�     NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�X`     NNNNNNNNNNNNNG�]�     G�^      G�^`     G�^�     G�_      G�_�     G�_�     G�`      G�`P     G�`�     G�`�     G�`�     G�a     G�a@     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNG�X      NNNNNNNNNNNNNG�]@     NNNNNNG�`P     G�`�     G�`�     G�`�     G�a     G�a@     G�ap     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�V�     G�W@     G�W�     G�X      G�X`     G�X�     NNNNNNNNNNG�\�     NNNNNNG�`�     G�`�     G�`�     G�a     G�a@     G�ap     G�a�     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�V�     G�V�     G�W@     G�W�     G�X      G�X`     NNNNNNNNNNG�\�     NNNNNNG�`�     G�`�     G�a     G�a@     G�ap     G�a�     G�a�     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�V      G�V�     G�V�     G�W@     G�W�     G�X      NNNNNNNNNNG�\      NNNNNNG�`�     G�a     G�a@     G�ap     G�a�     G�a�     G�b      NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�U�     G�V      G�V�     G�V�     G�W@     G�W�     G�X      G�X`     G�X�     G�Y      G�Y�     G�Y�     G�Z@     G�Z�     G�[      G�[`     G�[�     NNNNNNG�a     G�a@     G�ap     G�a�     G�a�     G�b      G�b0     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�U`     G�U�     G�V      G�V�     G�V�     G�W@     NNNNNNNNNNNNNNNNNG�a@     G�ap     G�a�     G�a�     G�b      G�b0     G�b`     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�U      G�U`     G�U�     G�V      G�V�     G�V�     NNNNNNNNNNNNNNNNNG�ap     G�a�     G�a�     G�b      G�b0     G�b`     G�b�     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�T�     G�U      G�U`     G�U�     G�V      G�V�     NNNNNNNNNNNNNNNNNG�a�     G�a�     G�b      G�b0     G�b`     G�b�     G�b�     NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�T@     G�T�     G�U      G�U`     G�U�     G�V      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�S�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�S�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�S      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�R�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNG�R`     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNG�P�     G�Q@     G�Q�     G�R      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�      G�      G��      G�      NNNNNNNNNNNNNNNNNNe]�(NNNNG�P�     NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�      G�      G��      G�       G��      NNNNNNNNNNNNNNNNNNe]�(NNNNG�P      NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�      G�      G�      G�      G��      G�      NNNNNNNNNNNNNNNNNNe]�(NNNNG�O�     G�N�     G�N      G�M@     G�L�     NNNNNNNNNNNNNNNNNNNNNNNNNNNG�"      G�      G�      G�      G�      G�      NNNNNNNNNNNNNNNNNNe]�(NNNNG�N�     G�N      G�M@     G�L�     G�K�     G�K      G�J@     G�I�     G�H�     G�H      G�G@     G�F�     G�E�     G�E      G�D@     G�C�     NNNNNNNNNNNNNNNNG�%      G�"      G�      G�      G�      G�      NNNNNNNNNNNNNNNNNNe]�(NNNNG�O�     G�N�     G�N      G�M@     G�L�     NNNNNNNNNNG�B�     G�B      G�A@     G�@�     G�?�     G�>      G�<�     G�;      G�9�     G�8      G�6�     G�5      G�3�     G�2      G�0�     G�.      G�+      G�(      G�%      G�"      G�      G�      G�      NNNNNNNNNNNNNNNNNNe]�(NNNNG�P      G�O�     G�N�     G�N      G�M@     NNNNNNNNNNNNNNNNNNNNNNNNNNNG�+      G�(      G�%      G�"      G�      G�"      NNNNNNNNNNNNNNNNNNe]�(NNNNG�P�     G�P      G�O�     G�N�     G�N      NNNNNNNNNNNNNNNNNNNNNNNNNNNG�.      G�+      G�(      G�%      G�"      G�%      NNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNG�0�     G�.      G�+      G�(      G�%      G�(      NNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej�{  ]�(j4,  j�-  jA.  ej�{  j�{  j�{  ]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKKKKK KK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K KKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKK K K K K K K K KKKKKKKKKKKKKKKKKKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K KKKKKKKK K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K eej�{  ]�(]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j.,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j<,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  jF,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j<,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  jV,  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j.,  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  jV,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  jF,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j.,  j�{  j�{  j�{  j�-  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j,  jV,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  jV,  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  e]�(j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  j�{  eej5|  j�+  j6|  j�,  j7|  ]�(j�+  j�+  j�+  j�+  j�+  ej9|  ]�j;|  ]�(K(K)ej=|  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKKKKNNNNNNNNNNNKKKKKKKKKKKKK K!K"K#K$K%K&NNNNNNNNNNNNNNNNNNNNNNe]�(NNNKKKKKNNNNNNNNNNNKNNNNNNNNNNK K!K"K#K$K%K&K'NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNKNNNNNNNNNNK!K"K#K$K%K&K'K(NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKK KNNNNNNNNNNNKNNNNNNNNNNK"K#K$K%K&K'K(K)NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNKNNNNNNNNNNNK$K%K&K'K(K)K*NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKKKKKKK	K
KKKKKNNNNNNNNNNNNK&K'K(K)K*K+NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNK(NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNK)NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNK	KKKKKNNNNNNNNNNNNNNNNNNNNNNNNNK*NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK+NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK,NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK-NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK	NNNNNNNNNNNNNNNNNNNNNNNNNNK.NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK
NNNNNNNNNNNNNNNNNNNNNNNNNNK/NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKKKKNNNNNNNNNNNNNNNNNNNNNNNK0NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK5NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNK,K-K.K/K0K1K2K3K4K5K6K7K8K9NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNK+NNNNNNK4K5K6K7K8K9K:NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNK*NNNNNNK5K6K7K8K9K:K;NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNK)NNNNNNK6K7K8K9K:K;K<NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNK(NNNNNNK7K8K9K:K;K<K=NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKKKKK K!K"K#K$K%K&K'NNNNNNK8K9K:K;K<K=K>NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNK9K:K;K<K=K>K?NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNK:K;K<K=K>K?K@NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNK;K<K=K>K?K@KANNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKK NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK!NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK"NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK#NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK$NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNK(K'K&K%NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKTKUKVKWNNNNNNNNNNNNNNNNNNe]�(NNNNK)NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKRKSKTKUKVNNNNNNNNNNNNNNNNNNe]�(NNNNK*NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKPKQKRKSKTKUNNNNNNNNNNNNNNNNNNe]�(NNNNK+K,K-K.K/NNNNNNNNNNNNNNNNNNNNNNNNNNNKOKPKQKRKSKTNNNNNNNNNNNNNNNNNNe]�(NNNNK,K-K.K/K0K1K2K3K4K5K6K7K8K9K:K;NNNNNNNNNNNNNNNNKNKOKPKQKRKSNNNNNNNNNNNNNNNNNNe]�(NNNNK-K.K/K0K1NNNNNNNNNNK<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQKRNNNNNNNNNNNNNNNNNNe]�(NNNNK.K/K0K1K2NNNNNNNNNNNNNNNNNNNNNNNNNNNKNKOKPKQKRKSNNNNNNNNNNNNNNNNNNe]�(NNNNK/K0K1K2K3NNNNNNNNNNNNNNNNNNNNNNNNNNNKOKPKQKRKSKTNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKPKQKRKSKTKUNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej�|  hj�|  ]�(]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNKKKKNNNNNNNNNNNKKKKKKKKKKKKKK K!K"K#K$K%NNNNNNNNNNNNNNNNNNNNNNe]�(NNNKKKKKNNNNNNNNNNNKNNNNNNNNNNKK K!K"K#K$K%K&NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKK KNNNNNNNNNNNKNNNNNNNNNNK K!K"K#K$K%K&K'NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKK KK NNNNNNNNNNNKNNNNNNNNNNK!K"K#K$K%K&K'K(NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKK KNNNNNNNNNNNKNNNNNNNNNNNK#K$K%K&K'K(K)NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKKKKKKKK	K
KKKKNNNNNNNNNNNNK%K&K'K(K)K*NNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNK'NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNK(NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNK)NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK*NNNN�~*      NNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK+NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK,NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNK-NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK	NNNNNNNNNNNNNNNNNNNNNNNNNNK.NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNK
KKKNNNNNNNNNNNNNNNNNNNNNNNK/NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK0NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK1NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK2NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK3NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNK4NNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNK+K,K-K.K/K0K1K2K3K4K5K6K7K8NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNKNNNNNNNNNNNNNK*NNNNNNK3K4K5K6K7K8K9NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNK)NNNNNNK4K5K6K7K8K9K:NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNK(NNNNNNK5K6K7K8K9K:K;NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNK'NNNNNNK6K7K8K9K:K;K<NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKKKKKK K!K"K#K$K%K&NNNNNNK7K8K9K:K;K<K=NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNK8K9K:K;K<K=K>NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNK9K:K;K<K=K>K?NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNK:K;K<K=K>K?K@NNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKKKKKKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNKNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK!NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK"NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNK#NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNK'K&K%K$NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKSKTKUKVNNNNNNNNNNNNNNNNNNe]�(NNNNK(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKQKRKSKTKUNNNNNNNNNNNNNNNNNNe]�(NNNNK)NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKOKPKQKRKSKTNNNNNNNNNNNNNNNNNNe]�(NNNNK*K+K,K-K.NNNNNNNNNNNNNNNNNNNNNNNNNNNKNKOKPKQKRKSNNNNNNNNNNNNNNNNNNe]�(NNNNK+K,K-K.K/K0K1K2K3K4K5K6K7K8K9K:NNNNNNNNNNNNNNNNKMKNKOKPKQKRNNNNNNNNNNNNNNNNNNe]�(NNNNK,K-K.K/K0NNNNNNNNNNK;K<K=K>K?K@KAKBKCKDKEKFKGKHKIKJKKKLKMKNKOKPKQNNNNNNNNNNNNNNNNNNe]�(NNNNK-K.K/K0K1NNNNNNNNNNNNNNNNNNNNNNNNNNNKMKNKOKPKQKRNNNNNNNNNNNNNNNNNNe]�(NNNNK.K/K0K1K2NNNNNNNNNNNNNNNNNNNNNNNNNNNKNKOKPKQKRKSNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNKOKPKQKRKSKTNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNe]�(NNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNNeej�|  jK�  j7,  �1B: Dark Crypt�j�|  j�|  jX}  ]�(]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKKK K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K KKKKKKKK K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K e]�(K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K K eej�}  Jv j�}  j�}  ubj]-  ej�|  j�|  j�|  h�cursor�Kub�width�K#�turn�M��xConst�Kj6|  j�,  �yConst�KF�height�K�MessageHandler�j�|  ub.